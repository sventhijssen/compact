// IWLS benchmark module "x1" printed on Wed May 29 16:25:46 2002
module x1(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2, b2, c2, d2, e2, f2, g2, h2, i2);
input
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  t,
  u,
  v,
  w,
  y,
  z,
  a0,
  b0,
  c0,
  d0,
  e0,
  f0,
  g0,
  h0,
  i0,
  j0,
  k0,
  l0,
  m0,
  n0,
  o0,
  p0,
  q0,
  r0,
  s0,
  t0,
  u0,
  v0,
  w0,
  x0,
  y0,
  z0;
output
  a1,
  a2,
  b1,
  b2,
  c1,
  c2,
  d1,
  d2,
  e1,
  e2,
  f1,
  f2,
  g1,
  g2,
  h1,
  h2,
  i1,
  i2,
  j1,
  k1,
  l1,
  m1,
  n1,
  o1,
  p1,
  q1,
  r1,
  s1,
  t1,
  u1,
  v1,
  w1,
  x1,
  y1,
  z1;
wire
  \[5] ,
  \[6] ,
  \[7] ,
  \[21] ,
  \[22] ,
  \[23] ,
  \[24] ,
  \[25] ,
  \[26] ,
  \[27] ,
  \[29] ,
  \[30] ,
  \[31] ,
  \[32] ,
  \[33] ,
  \[34] ,
  \[10] ,
  \[11] ,
  \[12] ,
  \[13] ,
  \[14] ,
  \[0] ,
  \[1] ,
  \[17] ,
  \[2] ,
  \[18] ,
  \[3] ,
  \[4] ;
assign
  \[5]  = (e0 & (p & (~m & (~h & (~a & o))))) | ((~i & (~q & q0)) | ((~i & (q0 & ~o)) | ((~q & (q0 & ~g)) | (q0 & (~o & ~g))))),
  \[6]  = (~s & (~d & (p0 & (~q & (~h & (~g & (~a & (~v & ~m)))))))) | ((~s & (~d & (p0 & (~h & (~g & (~a & (~v & (~p & ~m)))))))) | ((~s & (~d & (p0 & (~h & (~g & (~a & (~v & (~o & ~m)))))))) | ((~s & (p0 & (~q & (~h & (~g & (~c & (~a & (~v & ~m)))))))) | ((~s & (p0 & (~h & (~g & (~c & (~a & (~v & (~p & ~m)))))))) | ((~s & (p0 & (~h & (~g & (~c & (~a & (~v & (~o & ~m)))))))) | ((~d & (p0 & (~r & (~q & (~h & (~g & (~a & (~v & ~m)))))))) | ((~d & (p0 & (~r & (~h & (~g & (~a & (~v & (~p & ~m)))))))) | ((~d & (p0 & (~r & (~h & (~g & (~a & (~v & (~o & ~m)))))))) | ((p0 & (~r & (~q & (~h & (~g & (~c & (~a & (~v & ~m)))))))) | ((p0 & (~r & (~h & (~g & (~c & (~a & (~v & (~p & ~m)))))))) | ((p0 & (~r & (~h & (~g & (~c & (~a & (~v & (~o & ~m)))))))) | ((~s & (~i & (p0 & (~q & (~h & (g & ~a)))))) | ((~s & (~i & (p0 & (~q & (~h & (~a & v)))))) | ((~s & (~i & (p0 & (~h & (g & (~a & ~p)))))) | ((~s & (~i & (p0 & (~h & (g & (~a & ~o)))))) | ((~s & (~i & (p0 & (~h & (~a & (v & ~p)))))) | ((~s & (~i & (p0 & (~h & (~a & (v & ~o)))))) | ((~i & (p0 & (~r & (~q & (~h & (g & ~a)))))) | ((~i & (p0 & (~r & (~q & (~h & (~a & v)))))) | ((~i & (p0 & (~r & (~h & (g & (~a & ~p)))))) | ((~i & (p0 & (~r & (~h & (g & (~a & ~o)))))) | ((~i & (p0 & (~r & (~h & (~a & (v & ~p)))))) | ((~i & (p0 & (~r & (~h & (~a & (v & ~o)))))) | ((g & (d0 & (~v & (u & (p & (o & ~m)))))) | ((g & (d0 & (~v & (p & (o & (~m & e)))))) | ((d0 & (~v & (~u & (p & (o & (~m & ~e)))))) | ((v0 & o0) | (d0 & v)))))))))))))))))))))))))))),
  \[7]  = (e0 & (~o & (~w & (~u & (h & (~e & ~a)))))) | ((d0 & (~d & (~w & (~u & (h & (~e & ~a)))))) | ((p0 & (~w & (~u & (h & (~e & ~a))))) | (s0 & (~w & (~u & (h & (~e & ~a))))))),
  \[21]  = (~f & (g0 & (v & (~m & (~j & ~a))))) | ((~r & (k0 & (~v & (~m & (~j & ~a))))) | ((k0 & (v & (n & (~m & (~j & ~a))))) | (g0 & (~v & (~m & (~j & ~a)))))),
  \[22]  = (k0 & (s & r)) | (a0 & (s & r)),
  \[23]  = (r0 & ~j) | ((f0 & ~j) | ((g0 & ~j) | (h0 | z))),
  \[24]  = (~r0 & (~g0 & (~f0 & (~h0 & ~z)))) | (~h0 & (~z & j)),
  \[25]  = c0 | d0,
  \[26]  = r0 | f0,
  \[27]  = (p0 & (~w & (~v & (~u & (p & (o & (~m & (~g & (~e & ~a))))))))) | ((e0 & (~w & (~v & (~u & (p & (o & (~m & (~g & (~e & ~a))))))))) | ((p0 & (~w & (~v & (~u & (~p & (o & (~m & (~e & ~a)))))))) | (e0 & (~w & (~v & (~u & (~p & (o & (~m & (~e & ~a)))))))))),
  \[29]  = (~o & (q0 & (~v & (i & (g & ~a))))) | ((~p & (q0 & (~v & (i & (g & ~a))))) | ((q0 & (~v & (~q & (i & (g & ~a))))) | ((p0 & (~o & (i & (g & ~a)))) | ((p0 & (~p & (i & (g & ~a)))) | ((p0 & (~q & (i & (g & ~a)))) | ((p0 & (v & (i & ~a))) | (y | (z | (h0 | i0))))))))),
  a1 = \[0] ,
  a2 = \[26] ,
  b1 = \[1] ,
  b2 = \[27] ,
  c1 = \[2] ,
  c2 = h0,
  d1 = \[3] ,
  d2 = \[29] ,
  e1 = \[4] ,
  e2 = \[30] ,
  f1 = \[5] ,
  f2 = \[31] ,
  g1 = \[6] ,
  \[30]  = (q & (p & (o & (~p0 & (~i0 & (~h0 & (~z & ~y))))))) | ((q & (p & (o & (~v & (~i0 & (~h0 & (~z & ~y))))))) | ((~q0 & (~p0 & (~i0 & (~h0 & (~z & ~y))))) | ((~p0 & (v & (~i0 & (~h0 & (~z & ~y))))) | ((~p0 & (~g & (~i0 & (~h0 & (~z & ~y))))) | ((~v & (~g & (~i0 & (~h0 & (~z & ~y))))) | ((~i & (~i0 & (~h0 & (~z & ~y)))) | (~i0 & (~h0 & (~z & (~y & a)))))))))),
  g2 = \[32] ,
  h1 = \[7] ,
  \[31]  = (r & (~m & (l & (~j & (b & (~t & (~e0 & (d & (~x0 & (~s0 & (~r0 & (~p0 & (~m0 & ~f0))))))))))))) | ((r & (~m & (l & (~j & (b & (~t & (~e0 & (~x0 & (~s0 & (~r0 & (~p0 & (~m0 & (~f0 & ~d0))))))))))))) | ((r & (~m & (l & (~j & (b & (~t & (d & (~x0 & (~s0 & (~r0 & (~p0 & (~m0 & (~f0 & o))))))))))))) | ((r & (~m & (l & (~j & (b & (~t & (~x0 & (~s0 & (~r0 & (~p0 & (~m0 & (~f0 & (~d0 & o))))))))))))) | ((r & (~m & (l & (~j & (b & (~e0 & (d & (~x0 & (~s0 & (~r0 & (~p0 & (~m0 & (~i0 & ~f0))))))))))))) | ((r & (~m & (l & (~j & (b & (~e0 & (~x0 & (~s0 & (~r0 & (~p0 & (~m0 & (~i0 & (~f0 & ~d0))))))))))))) | ((r & (~m & (l & (~j & (b & (d & (~x0 & (~s0 & (~r0 & (~p0 & (~m0 & (~i0 & (~f0 & o))))))))))))) | ((r & (~m & (l & (~j & (b & (~x0 & (~s0 & (~r0 & (~p0 & (~m0 & (~i0 & (~f0 & (~d0 & o))))))))))))) | ((z0 & (l & (b & (~t & (~e0 & (d & (~x0 & (~s0 & (~r0 & (~p0 & (~m0 & ~f0))))))))))) | ((z0 & (l & (b & (~t & (~e0 & (~x0 & (~s0 & (~r0 & (~p0 & (~m0 & (~f0 & ~d0))))))))))) | ((z0 & (l & (b & (~t & (d & (~x0 & (~s0 & (~r0 & (~p0 & (~m0 & (~f0 & o))))))))))) | ((z0 & (l & (b & (~t & (~x0 & (~s0 & (~r0 & (~p0 & (~m0 & (~f0 & (~d0 & o))))))))))) | ((z0 & (l & (b & (~e0 & (d & (~x0 & (~s0 & (~r0 & (~p0 & (~m0 & (~i0 & ~f0))))))))))) | ((z0 & (l & (b & (~e0 & (~x0 & (~s0 & (~r0 & (~p0 & (~m0 & (~i0 & (~f0 & ~d0))))))))))) | ((z0 & (l & (b & (d & (~x0 & (~s0 & (~r0 & (~p0 & (~m0 & (~i0 & (~f0 & o))))))))))) | ((z0 & (l & (b & (~x0 & (~s0 & (~r0 & (~p0 & (~m0 & (~i0 & (~f0 & (~d0 & o))))))))))) | ((r & (~m & (l & (~j & (b & (~h & (~x0 & (~r0 & (~m0 & ~f0))))))))) | ((~t & (~e0 & (d & (~x0 & (~s0 & (~r0 & (~p0 & (~m0 & (~f0 & ~a0))))))))) | ((~t & (~e0 & (~x0 & (~s0 & (~r0 & (~p0 & (~m0 & (~f0 & (~d0 & ~a0))))))))) | ((~t & (d & (~x0 & (~s0 & (~r0 & (~p0 & (~m0 & (~f0 & (~a0 & o))))))))) | ((~t & (~x0 & (~s0 & (~r0 & (~p0 & (~m0 & (~f0 & (~d0 & (~a0 & o))))))))) | ((~e0 & (d & (~x0 & (~s0 & (~r0 & (~p0 & (~m0 & (~i0 & (~f0 & ~a0))))))))) | ((~e0 & (~x0 & (~s0 & (~r0 & (~p0 & (~m0 & (~i0 & (~f0 & (~d0 & ~a0))))))))) | ((d & (~x0 & (~s0 & (~r0 & (~p0 & (~m0 & (~i0 & (~f0 & (~a0 & o))))))))) | ((~x0 & (~s0 & (~r0 & (~p0 & (~m0 & (~i0 & (~f0 & (~d0 & (~a0 & o))))))))) | ((z0 & (l & (b & (~h & (~x0 & (~r0 & (~m0 & ~f0))))))) | (~h & (~x0 & (~r0 & (~m0 & (~f0 & ~a0)))))))))))))))))))))))))))))),
  h2 = \[33] ,
  i1 = m0,
  \[32]  = (j & (~z0 & (a0 & b))) | ((m & (~z0 & (a0 & b))) | ((~z0 & (~r & (a0 & b))) | ((d0 & (~d & h)) | ((e0 & (~o & h)) | ((i0 & (t & h)) | ((a0 & (~l & b)) | ((s0 & h) | ((p0 & h) | ((a0 & ~b) | (m0 | (x0 | (r0 | f0)))))))))))),
  i2 = \[34] ,
  j1 = n0,
  \[33]  = (~k0 & (~g0 & (~a0 & (~i0 & (~h0 & (~c0 & (~b0 & (~z & (~y & (h & ~d)))))))))) | ((~k0 & (~g0 & (~a0 & (~h0 & (~c0 & (~b0 & (~z & (~y & (~i & (h & ~d)))))))))) | ((~k0 & (~a0 & (~i0 & (~c & (~h0 & (~c0 & (~b0 & (~z & (~y & (h & ~d)))))))))) | ((~k0 & (~a0 & (~i0 & (~h0 & (~c0 & (~b0 & (~z & (~y & (~j & (h & ~d)))))))))) | ((~k0 & (~a0 & (~c & (~h0 & (~c0 & (~b0 & (~z & (~y & (~i & (h & ~d)))))))))) | ((~k0 & (~a0 & (~h0 & (~c0 & (~b0 & (~z & (~y & (~j & (~i & (h & ~d)))))))))) | ((~v & (~g0 & (~a0 & (~i0 & (~h0 & (~c0 & (~b0 & (~z & (~y & (h & ~d)))))))))) | ((~v & (~g0 & (~a0 & (~h0 & (~c0 & (~b0 & (~z & (~y & (~i & (h & ~d)))))))))) | ((~v & (~a0 & (~i0 & (~c & (~h0 & (~c0 & (~b0 & (~z & (~y & (h & ~d)))))))))) | ((~v & (~a0 & (~c & (~h0 & (~c0 & (~b0 & (~z & (~y & (~i & (h & ~d)))))))))) | ((~g0 & (~a0 & (~i0 & (~h0 & (~c0 & (~b0 & (~z & (~y & (j & (h & ~d)))))))))) | ((~g0 & (~a0 & (~h0 & (~c0 & (~b0 & (~z & (~y & (j & (~i & (h & ~d)))))))))) | ((~a0 & (~i0 & (~c & (~h0 & (~c0 & (~b0 & (~z & (~y & (j & (h & ~d)))))))))) | ((~a0 & (~c & (~h0 & (~c0 & (~b0 & (~z & (~y & (j & (~i & (h & ~d)))))))))) | ((~k0 & (~g0 & (~a0 & (~i0 & (~d0 & (~h0 & (~c0 & (~b0 & (~z & ~y))))))))) | ((~k0 & (~g0 & (~a0 & (~d0 & (~h0 & (~c0 & (~b0 & (~z & (~y & ~i))))))))) | ((~k0 & (~a0 & (~i0 & (~d0 & (~c & (~h0 & (~c0 & (~b0 & (~z & ~y))))))))) | ((~k0 & (~a0 & (~i0 & (~d0 & (~h0 & (~c0 & (~b0 & (~z & (~y & ~j))))))))) | ((~k0 & (~a0 & (~d0 & (~c & (~h0 & (~c0 & (~b0 & (~z & (~y & ~i))))))))) | ((~k0 & (~a0 & (~d0 & (~h0 & (~c0 & (~b0 & (~z & (~y & (~j & ~i))))))))) | ((n & (~g0 & (~i0 & (~h0 & (~c0 & (~b0 & (~z & (~y & (h & ~d))))))))) | ((n & (~g0 & (~h0 & (~c0 & (~b0 & (~z & (~y & (~i & (h & ~d))))))))) | ((n & (~i0 & (~c & (~h0 & (~c0 & (~b0 & (~z & (~y & (h & ~d))))))))) | ((n & (~i0 & (~h0 & (~c0 & (~b0 & (~z & (~y & (~j & (h & ~d))))))))) | ((n & (~c & (~h0 & (~c0 & (~b0 & (~z & (~y & (~i & (h & ~d))))))))) | ((n & (~h0 & (~c0 & (~b0 & (~z & (~y & (~j & (~i & (h & ~d))))))))) | ((m & (~g0 & (~i0 & (~h0 & (~c0 & (~b0 & (~z & (~y & (h & ~d))))))))) | ((m & (~g0 & (~h0 & (~c0 & (~b0 & (~z & (~y & (~i & (h & ~d))))))))) | ((m & (~i0 & (~c & (~h0 & (~c0 & (~b0 & (~z & (~y & (h & ~d))))))))) | ((m & (~i0 & (~h0 & (~c0 & (~b0 & (~z & (~y & (~j & (h & ~d))))))))) | ((m & (~c & (~h0 & (~c0 & (~b0 & (~z & (~y & (~i & (h & ~d))))))))) | ((m & (~h0 & (~c0 & (~b0 & (~z & (~y & (~j & (~i & (h & ~d))))))))) | ((a & (~g0 & (~i0 & (~h0 & (~c0 & (~b0 & (~z & (~y & (h & ~d))))))))) | ((a & (~g0 & (~h0 & (~c0 & (~b0 & (~z & (~y & (~i & (h & ~d))))))))) | ((a & (~i0 & (~c & (~h0 & (~c0 & (~b0 & (~z & (~y & (h & ~d))))))))) | ((a & (~i0 & (~h0 & (~c0 & (~b0 & (~z & (~y & (~j & (h & ~d))))))))) | ((a & (~c & (~h0 & (~c0 & (~b0 & (~z & (~y & (~i & (h & ~d))))))))) | ((a & (~h0 & (~c0 & (~b0 & (~z & (~y & (~j & (~i & (h & ~d))))))))) | ((~v & (~g0 & (~a0 & (~i0 & (~d0 & (~h0 & (~c0 & (~b0 & (~z & ~y))))))))) | ((~v & (~g0 & (~a0 & (~d0 & (~h0 & (~c0 & (~b0 & (~z & (~y & ~i))))))))) | ((~v & (~a0 & (~i0 & (~d0 & (~c & (~h0 & (~c0 & (~b0 & (~z & ~y))))))))) | ((~v & (~a0 & (~d0 & (~c & (~h0 & (~c0 & (~b0 & (~z & (~y & ~i))))))))) | ((~v & (~i0 & (~h0 & (~c0 & (~b0 & (~z & (~y & (~j & (h & ~d))))))))) | ((~v & (~h0 & (~c0 & (~b0 & (~z & (~y & (~j & (~i & (h & ~d))))))))) | ((~g0 & (~a0 & (~i0 & (~d0 & (~h0 & (~c0 & (~b0 & (~z & (~y & j))))))))) | ((~g0 & (~a0 & (~d0 & (~h0 & (~c0 & (~b0 & (~z & (~y & (j & ~i))))))))) | ((~g0 & (~i0 & (~b & (~h0 & (~c0 & (~b0 & (~z & (~y & (h & ~d))))))))) | ((~g0 & (~i0 & (~h0 & (~c0 & (~b0 & (~z & (~y & (~l & (h & ~d))))))))) | ((~g0 & (~b & (~h0 & (~c0 & (~b0 & (~z & (~y & (~i & (h & ~d))))))))) | ((~g0 & (~h0 & (~c0 & (~b0 & (~z & (~y & (~l & (~i & (h & ~d))))))))) | ((~a0 & (~i0 & (~d0 & (~c & (~h0 & (~c0 & (~b0 & (~z & (~y & j))))))))) | ((~a0 & (~d0 & (~c & (~h0 & (~c0 & (~b0 & (~z & (~y & (j & ~i))))))))) | ((~i0 & (~c & (~b & (~h0 & (~c0 & (~b0 & (~z & (~y & (h & ~d))))))))) | ((~i0 & (~c & (~h0 & (~c0 & (~b0 & (~z & (~y & (~l & (h & ~d))))))))) | ((~i0 & (~b & (~h0 & (~c0 & (~b0 & (~z & (~y & (~j & (h & ~d))))))))) | ((~i0 & (~h0 & (~c0 & (~b0 & (~z & (~y & (~l & (~j & (h & ~d))))))))) | ((~c & (~b & (~h0 & (~c0 & (~b0 & (~z & (~y & (~i & (h & ~d))))))))) | ((~c & (~h0 & (~c0 & (~b0 & (~z & (~y & (~l & (~i & (h & ~d))))))))) | ((~b & (~h0 & (~c0 & (~b0 & (~z & (~y & (~j & (~i & (h & ~d))))))))) | ((~h0 & (~c0 & (~b0 & (~z & (~y & (~l & (~j & (~i & (h & ~d))))))))) | ((n & (~g0 & (~i0 & (~d0 & (~h0 & (~c0 & (~b0 & (~z & ~y)))))))) | ((n & (~g0 & (~d0 & (~h0 & (~c0 & (~b0 & (~z & (~y & ~i)))))))) | ((n & (~i0 & (~d0 & (~c & (~h0 & (~c0 & (~b0 & (~z & ~y)))))))) | ((n & (~i0 & (~d0 & (~h0 & (~c0 & (~b0 & (~z & (~y & ~j)))))))) | ((n & (~d0 & (~c & (~h0 & (~c0 & (~b0 & (~z & (~y & ~i)))))))) | ((n & (~d0 & (~h0 & (~c0 & (~b0 & (~z & (~y & (~j & ~i)))))))) | ((m & (~g0 & (~i0 & (~d0 & (~h0 & (~c0 & (~b0 & (~z & ~y)))))))) | ((m & (~g0 & (~d0 & (~h0 & (~c0 & (~b0 & (~z & (~y & ~i)))))))) | ((m & (~i0 & (~d0 & (~c & (~h0 & (~c0 & (~b0 & (~z & ~y)))))))) | ((m & (~i0 & (~d0 & (~h0 & (~c0 & (~b0 & (~z & (~y & ~j)))))))) | ((m & (~d0 & (~c & (~h0 & (~c0 & (~b0 & (~z & (~y & ~i)))))))) | ((m & (~d0 & (~h0 & (~c0 & (~b0 & (~z & (~y & (~j & ~i)))))))) | ((a & (~g0 & (~i0 & (~d0 & (~h0 & (~c0 & (~b0 & (~z & ~y)))))))) | ((a & (~g0 & (~d0 & (~h0 & (~c0 & (~b0 & (~z & (~y & ~i)))))))) | ((a & (~i0 & (~d0 & (~c & (~h0 & (~c0 & (~b0 & (~z & ~y)))))))) | ((a & (~i0 & (~d0 & (~h0 & (~c0 & (~b0 & (~z & (~y & ~j)))))))) | ((a & (~d0 & (~c & (~h0 & (~c0 & (~b0 & (~z & (~y & ~i)))))))) | ((a & (~d0 & (~h0 & (~c0 & (~b0 & (~z & (~y & (~j & ~i)))))))) | ((~v & (~i0 & (~d0 & (~h0 & (~c0 & (~b0 & (~z & (~y & ~j)))))))) | ((~v & (~d0 & (~h0 & (~c0 & (~b0 & (~z & (~y & (~j & ~i)))))))) | ((~g0 & (~i0 & (~d0 & (~b & (~h0 & (~c0 & (~b0 & (~z & ~y)))))))) | ((~g0 & (~i0 & (~d0 & (~h0 & (~c0 & (~b0 & (~z & (~y & ~l)))))))) | ((~g0 & (~d0 & (~b & (~h0 & (~c0 & (~b0 & (~z & (~y & ~i)))))))) | ((~g0 & (~d0 & (~h0 & (~c0 & (~b0 & (~z & (~y & (~l & ~i)))))))) | ((~i0 & (~d0 & (~c & (~b & (~h0 & (~c0 & (~b0 & (~z & ~y)))))))) | ((~i0 & (~d0 & (~c & (~h0 & (~c0 & (~b0 & (~z & (~y & ~l)))))))) | ((~i0 & (~d0 & (~b & (~h0 & (~c0 & (~b0 & (~z & (~y & ~j)))))))) | ((~i0 & (~d0 & (~h0 & (~c0 & (~b0 & (~z & (~y & (~l & ~j)))))))) | ((~d0 & (~c & (~b & (~h0 & (~c0 & (~b0 & (~z & (~y & ~i)))))))) | ((~d0 & (~c & (~h0 & (~c0 & (~b0 & (~z & (~y & (~l & ~i)))))))) | ((~d0 & (~b & (~h0 & (~c0 & (~b0 & (~z & (~y & (~j & ~i)))))))) | (~d0 & (~h0 & (~c0 & (~b0 & (~z & (~y & (~l & (~j & ~i)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))),
  k1 = \[10] ,
  \[34]  = (k0 & (v & (~n & (~m & (l & (b & (~a & (g0 & c)))))))) | ((k0 & (v & (~n & (~m & (l & (b & (~a & ~j))))))) | ((a0 & (v & (~n & (~m & (l & (b & ~a)))))) | ((a0 & (~n & (~m & (l & (b & (~a & j)))))) | ((g0 & (j & c)) | ((d & d0) | ((d0 & ~h) | ((i0 & i) | (y | (b0 | (c0 | (h0 | z))))))))))),
  l1 = \[11] ,
  m1 = \[12] ,
  n1 = \[13] ,
  o1 = \[14] ,
  p1 = y,
  q1 = z,
  \[10]  = (d0 & (w & (~v & d))) | ((~j & (a & g0)) | ((i0 & (t & a)) | ((l0 & (s & r)) | ((s & (r & p0)) | ((b0 & (~v & m)) | ((c0 & (~v & m)) | ((p0 & (~v & m)) | ((d0 & (~v & m)) | ((j0 & a) | ((a0 & a) | ((a & s0) | ((a & q0) | ((a & k0) | ((a & p0) | ((a & d0) | ((a & h0) | ((a & e0) | ((s0 & m) | ((q0 & m) | ((k0 & m) | ((r0 & b) | ((h0 & m) | ((g0 & m) | (e0 & m)))))))))))))))))))))))),
  r1 = \[17] ,
  \[11]  = (~v & (p & (o & (~g & (~d & (~a & (e & (d0 & ~h)))))))) | ((~v & (p & (o & (~g & (~d & (~a & (d0 & (u & ~h)))))))) | ((~v & (~p & (o & (d & (~a & (e & (d0 & ~h))))))) | ((~v & (~p & (o & (d & (~a & (d0 & (u & ~h))))))) | ((e0 & (~v & (~p & (o & (~a & (e & ~h)))))) | ((e0 & (~v & (~p & (o & (~a & (u & ~h)))))) | ((~v & (~g & (d & (~a & (e & (d0 & ~h)))))) | ((~v & (~g & (d & (~a & (d0 & (u & ~h)))))) | ((e0 & (~v & (~g & (~a & (e & ~h))))) | ((e0 & (~v & (~g & (~a & (u & ~h))))) | ((q0 & (q & (p & o))) | ((p0 & (q & (p & o))) | ((a0 & (k & b)) | ((e0 & (e & h)) | ((e0 & (u & h)) | ((e & (d0 & h)) | ((d0 & (u & h)) | ((f0 & b) | ((w & h0) | ((h0 & e) | (h0 & u)))))))))))))))))))),
  s1 = \[18] ,
  \[12]  = (d0 & (~w & (~v & (~u & (~p & (o & (~m & (~e & (d & ~a))))))))) | (h0 & j),
  t1 = x0,
  \[13]  = (p0 & (d & (~g & (~w & (~u & (~e & (~m & (c & (~v & ~a))))))))) | ((q0 & (~q & (~g & (~w & (~u & (p & (o & (~e & (~m & ~a))))))))) | ((e0 & (~w & (~u & (~p & (o & (~e & (~m & ~a))))))) | ((w0 & (o0 & (~w & (~u & (~e & (~m & ~a)))))) | ((s0 & (~w & (~u & (~e & (~m & (~h & ~a)))))) | ((h0 & (~w & (~u & (~e & (~m & (~j & ~a)))))) | ((~m & (~h & (~c & (g0 & (j & ~a))))) | (g0 & (v & (~j & (f & ~a)))))))))),
  u1 = y0,
  \[14]  = (~o & (q0 & (g & (~v & (i & ~a))))) | ((~o & (g & (p0 & (~v & (i & ~a))))) | ((~p & (q0 & (g & (~v & (i & ~a))))) | ((~p & (g & (p0 & (~v & (i & ~a))))) | ((q0 & (~q & (g & (~v & (i & ~a))))) | ((~q & (g & (p0 & (~v & (i & ~a))))) | ((p0 & (v & (i & ~a))) | (i0 & (i & (~h & ~a))))))))),
  v1 = \[21] ,
  \[0]  = (a0 & (~v & (~r & ~j))) | ((r0 & ~b) | ((f0 & ~b) | ((~b & a0) | ((~l & a0) | ((m & a0) | (n & a0)))))),
  w1 = \[22] ,
  \[1]  = (a0 & (l & (~k & (v & (~n & (~m & (~j & (b & ~a)))))))) | ((a0 & (l & (~k & (~n & (~m & (j & (b & ~a))))))) | ((k0 & (v & (~n & (~m & (~j & (b & ~a)))))) | ((g0 & (~w & (c & j))) | (t0 & o0)))),
  x1 = \[23] ,
  \[17]  = (a0 & (l & (~k & (~v & (~s & (r & (~m & (~j & (b & ~a))))))))) | ((k0 & (~v & (~s & (r & (~m & (~j & (b & ~a))))))) | ((~t & (i0 & (~i & (~h & a)))) | ((i0 & (~i & (~h & ~a))) | (j0 & ~a)))),
  \[2]  = (~m & (b0 & ~v)) | (b0 & v),
  y1 = \[24] ,
  \[18]  = i0 & (t & h),
  \[3]  = (~o & (d0 & (~h & (~d & (~a & (~m & ~v)))))) | ((d0 & (~p & (~h & (~d & (~a & (~m & ~v)))))) | ((~m & (c0 & ~v)) | (c0 & v))),
  z1 = \[25] ,
  \[4]  = (~w & (~e & (d0 & (~u & (~o & (~m & d)))))) | ((e & (d0 & (~o & (~m & (g & d))))) | ((d0 & (u & (~o & (~m & (g & d))))) | ((e0 & (~h & (~a & (~o & ~m)))) | (u0 & o0))));
endmodule

