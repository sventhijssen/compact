// IWLS benchmark module "lal" printed on Wed May 29 16:09:11 2002
module lal(a, b, c, d, e, f, g, h, j, k, l, m, n, o, p, q, r, s, t, u, v, w, \x , y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0);
input
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  t,
  u,
  v,
  w,
  \x ,
  y,
  z,
  a0;
output
  b0,
  c0,
  d0,
  e0,
  f0,
  g0,
  h0,
  i0,
  j0,
  k0,
  l0,
  m0,
  n0,
  o0,
  p0,
  q0,
  r0,
  s0,
  t0;
wire
  \[5] ,
  \[6] ,
  \[7] ,
  \[8] ,
  \[9] ,
  a2,
  a3,
  a4,
  b2,
  b3,
  c2,
  c3,
  d2,
  d3,
  d4,
  e3,
  f2,
  f3,
  f4,
  g2,
  g3,
  h2,
  i2,
  i3,
  j3,
  k2,
  k3,
  k4,
  l2,
  l3,
  m2,
  m3,
  n1,
  n2,
  n3,
  o2,
  o3,
  p2,
  p3,
  q1,
  \[10] ,
  r2,
  \[11] ,
  r3,
  s2,
  \[12] ,
  s3,
  t2,
  \[13] ,
  t3,
  u2,
  \[14] ,
  u3,
  v2,
  \[15] ,
  v3,
  \[0] ,
  w2,
  \[16] ,
  w3,
  \[1] ,
  x1,
  x2,
  \[17] ,
  x3,
  y1,
  \[18] ,
  \[3] ,
  z2,
  \[4] ;
assign
  \[5]  = ~j & ~o,
  \[6]  = ~j & p,
  \[7]  = ~k4,
  \[8]  = (~t3 & (~u3 & w)) | ~v3,
  \[9]  = ~n1 & ~q,
  a2 = s & (t & u),
  a3 = (~b3 & (~q & ~e)) | (~b3 & (~q & ~f)),
  a4 = (d & ~n) | ((c & ~m) | ~d4),
  b0 = \[0] ,
  b2 = (~c2 & (~q & ~e)) | (~c2 & (~q & ~f)),
  b3 = ~c3 & (~y & ~z),
  c0 = \[1] ,
  c2 = ~d2 & ~v,
  c3 = ~e3 | (~d3 | ~s),
  d0 = r,
  d2 = ~s | (~t | ~u),
  d3 = t & u,
  d4 = (~f4 & a) | (~f4 & ~k),
  e0 = \[3] ,
  e3 = ~v & (~w & ~\x ),
  f0 = \[4] ,
  f2 = ~i2 & (s & t),
  f3 = ~t | (~u | v),
  f4 = (n & ~d) | ((m & ~c) | (l & ~b)),
  g0 = \[5] ,
  g2 = (~h2 & (~q & ~e)) | (~h2 & (~q & ~f)),
  g3 = w | (\x  | y),
  h0 = \[6] ,
  h2 = ~d2 & (~v & ~w),
  i0 = \[7] ,
  i2 = ~u | v,
  i3 = ~p3 & (~p2 & ~o3),
  j0 = \[8] ,
  j3 = (~k3 & (~q & ~e)) | (~k3 & (~q & ~f)),
  k0 = \[9] ,
  k2 = ~p2 & (s & t),
  k3 = ~l3 & (~z & ~a0),
  k4 = g & ~j,
  l0 = \[10] ,
  l2 = (~m2 & (~q & ~e)) | (~m2 & (~q & ~f)),
  l3 = ~n3 | (~m3 | ~s),
  m0 = \[11] ,
  m2 = ~n2 & (~w & ~\x ),
  m3 = t & (u & ~v),
  n0 = \[12] ,
  n1 = ~e | (~f | h),
  n2 = ~o2 | (~s | ~t),
  n3 = ~w & (~\x  & ~y),
  o0 = \[13] ,
  o2 = u & ~v,
  o3 = ~s | ~t,
  p0 = \[14] ,
  p2 = ~u | (v | w),
  p3 = \x  | (y | z),
  q0 = \[15] ,
  q1 = (f & e) | (q | h),
  \[10]  = ~q1 & ~s,
  r0 = \[16] ,
  r2 = ~x2 & (~w2 & s),
  \[11]  = (~q1 & (~t & s)) | (~q1 & (t & ~s)),
  r3 = ~t3 & (w & \x ),
  s0 = \[17] ,
  s2 = (~t2 & (~q & ~e)) | (~t2 & (~q & ~f)),
  \[12]  = (~x1 & (t & s)) | (~x1 & u),
  s3 = (~h & (~f & a0)) | ((~h & (~f & z)) | ((~h & (~e & a0)) | (~h & (~e & z)))),
  t0 = \[18] ,
  t2 = ~u2 & (~\x  & ~y),
  \[13]  = (~a2 & v) | (~b2 | h),
  t3 = (~v & u) | ((~v & t) | (~v & s)),
  u2 = ~v2 | (~s | ~t),
  \[14]  = (~f2 & w) | (~g2 | h),
  u3 = ~\x  | ~z,
  v2 = u & (~v & ~w),
  \[15]  = (~k2 & \x ) | (~l2 | h),
  v3 = (~a0 & ~z) | (~a0 & ~y),
  \[0]  = j & ~r,
  w2 = ~t | ~u,
  \[16]  = (~r2 & y) | (~s2 | h),
  w3 = (~t3 & (~u3 & w)) | ~v3,
  \[1]  = (~r3 & (~y & ~a0)) | ~s3,
  x1 = (s & (t & u)) | ~y1,
  x2 = v | (w | \x ),
  \[17]  = (~z2 & z) | (~a3 | h),
  x3 = (~a4 & (~b & ~a)) | ((~a4 & (~b & k)) | ((~a4 & (l & ~a)) | (~a4 & (l & k)))),
  y1 = (~q & (~h & ~f)) | (~q & (~h & ~e)),
  \[18]  = (~i3 & a0) | (~j3 | h),
  \[3]  = ~w3,
  z2 = ~g3 & (~f3 & s),
  \[4]  = ~x3 & ~j;
endmodule

