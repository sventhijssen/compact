module s27(VDD,CK,G0,G1,G17,G2,G3);
input VDD,CK,G0,G1,G2,G3;
output G17;

  wire G5,G10,G6,G11,G7,G13,G14,G8,G15,G12,G16,G9;

  FD1 DFF_0(CK,G5,G10);
  FD1 DFF_1(CK,G6,G11);
  FD1 DFF_2(CK,G7,G13);
  IV  NOT_0(G14,G0);
  IV  NOT_1(G17,G11);
  AN2 AND2_0(G8,G14,G6);
  OR2 OR2_0(G15,G12,G8);
  OR2 OR2_1(G16,G3,G8);
  ND2 NAND2_0(G9,G16,G15);
  NR2 NOR2_0(G10,G14,G11);
  NR2 NOR2_1(G11,G5,G9);
  NR2 NOR2_2(G12,G1,G7);
  NR2 NOR2_3(G13,G2,G12);

endmodule
