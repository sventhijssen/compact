// IWLS benchmark module "c8" printed on Wed May 29 16:07:19 2002
module c8(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, u, v, w, \x , y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0);
input
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  u,
  v,
  w,
  \x ,
  y,
  z,
  a0,
  b0,
  c0;
output
  g0,
  h0,
  i0,
  j0,
  k0,
  l0,
  m0,
  n0,
  o0,
  p0,
  q0,
  r0,
  s0,
  t0,
  u0,
  d0,
  e0,
  f0;
wire
  \[26] ,
  h2,
  \[27] ,
  \[10] ,
  \[11] ,
  \[12] ,
  n2,
  \[13] ,
  \[14] ,
  \[0] ,
  \[15] ,
  \[1] ,
  \[16] ,
  \[2] ,
  \[17] ,
  \[3] ,
  \[18] ,
  t2,
  \[4] ,
  \[19] ,
  \[5] ,
  v1,
  \[6] ,
  \[7] ,
  \[9] ,
  z1,
  z2,
  \[20] ,
  \[21] ,
  \[22] ,
  d2,
  \[23] ,
  \[24] ,
  \[25] ;
assign
  g0 = \[3] ,
  \[26]  = \[24]  | w,
  h0 = \[4] ,
  h2 = (\[23]  & ~e) | (\[22]  & ~m),
  \[27]  = v | ~q,
  i0 = \[5] ,
  j0 = \[6] ,
  k0 = \[7] ,
  \[10]  = (\[27]  & ~v1) | (~\[20]  & ~v1),
  l0 = c0,
  \[11]  = (\[24]  & (~z1 & w)) | ((~\[26]  & ~z1) | (~z1 & ~q)),
  m0 = \[9] ,
  \[12]  = (\[26]  & (~d2 & \x )) | ((~\[18]  & ~d2) | (~d2 & ~q)),
  n0 = \[10] ,
  n2 = (\[23]  & ~f) | (\[22]  & ~n),
  \[13]  = (\[18]  & (~h2 & y)) | ((~\[19]  & ~h2) | (~h2 & ~q)),
  o0 = \[11] ,
  \[14]  = (\[19]  & (~n2 & z)) | ((~\[21]  & ~n2) | (~n2 & ~q)),
  p0 = \[12] ,
  \[0]  = (~c0 & ~u) | (c0 & ~i),
  \[15]  = (\[21]  & (~t2 & a0)) | ((~\[25]  & ~t2) | (~t2 & ~q)),
  q0 = \[13] ,
  \[1]  = (~c0 & ~v) | (c0 & ~j),
  \[16]  = (~\[25]  & (~z2 & ~b0)) | ((\[25]  & (~z2 & b0)) | (~z2 & ~q)),
  r0 = \[14] ,
  \[2]  = (~c0 & ~w) | (c0 & ~k),
  \[17]  = (~\[27]  & (~b0 & (~a0 & (~z & (~y & (~\x  & (~w & (u & ~r)))))))) | (c0 & (r & q)),
  s0 = \[15] ,
  \[3]  = (~c0 & ~\x ) | (c0 & ~l),
  \[18]  = \[20]  | (\x  | (w | v)),
  t0 = \[16] ,
  t2 = (\[23]  & ~g) | (\[22]  & ~o),
  \[4]  = (~c0 & ~y) | (c0 & ~m),
  \[19]  = \[18]  | y,
  u0 = \[17] ,
  \[5]  = (~c0 & ~z) | (c0 & ~n),
  v1 = (~\[20]  & (v & q)) | ((\[23]  & ~b) | (\[22]  & ~j)),
  \[6]  = (~c0 & ~a0) | (c0 & ~o),
  \[7]  = (~c0 & ~b0) | (c0 & ~p),
  \[9]  = (u & (r & q)) | ((\[23]  & a) | ((\[22]  & i) | (~\[20]  & q))),
  z1 = (\[23]  & ~c) | (\[22]  & ~k),
  z2 = (\[23]  & ~h) | (\[22]  & ~p),
  \[20]  = u | r,
  \[21]  = \[19]  | z,
  \[22]  = ~s & ~q,
  d0 = \[0] ,
  d2 = (\[23]  & ~d) | (\[22]  & ~l),
  \[23]  = s & ~q,
  e0 = \[1] ,
  \[24]  = \[20]  | v,
  f0 = \[2] ,
  \[25]  = \[21]  | a0;
endmodule

