// C432
module foobar(k0, l0, m0, n0, o0, p0, q0, a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0);
input a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0;
output k0, l0, m0, n0, o0, p0, q0;
not(k0, r2);
not(l0, f4);
not(m0, r5);
not(t_0, q6);
not(t_1, l6);
and(n0, t_0, t_1);
not(t_2, g6);
not(t_3, u6);
not(t_4, i6);
not(t_5, j6);
or(o0, t_2, t_3, t_4, t_5);
not(t_6, t6);
not(t_7, s6);
not(t_8, i6);
not(t_9, j6);
or(p0, t_6, t_7, t_8, t_9);
not(t_10, r6);
not(t_11, s6);
not(t_12, u6);
not(t_13, j6);
or(q0, t_10, t_11, t_12, t_13);
not(y0, h0);
not(z0, f0);
not(a1, d0);
not(b1, b0);
not(c1, z);
not(d1, x);
not(e1, v);
not(f1, t);
not(g1, r);
not(h1, p);
not(i1, n);
not(j1, l);
not(k1, j);
not(l1, h);
not(m1, f);
not(n1, d);
not(o1, b);
not(p1, a);
not(t_14, j0);
not(t_15, y0);
and(q1, t_14, t_15);
not(t_16, i0);
not(t_17, y0);
and(r1, t_16, t_17);
not(t_18, h0);
not(t_19, z0);
or(s1, t_18, t_19);
not(t_20, g0);
not(t_21, a1);
and(t1, t_20, t_21);
not(t_22, e0);
not(t_23, a1);
and(u1, t_22, t_23);
not(t_24, d0);
not(t_25, b1);
or(v1, t_24, t_25);
not(t_26, c0);
not(t_27, c1);
and(w1, t_26, t_27);
not(t_28, a0);
not(t_29, c1);
and(x1, t_28, t_29);
not(t_30, z);
not(t_31, d1);
or(y1, t_30, t_31);
not(t_32, y);
not(t_33, e1);
and(z1, t_32, t_33);
not(t_34, w);
not(t_35, e1);
and(a2, t_34, t_35);
not(t_36, v);
not(t_37, f1);
or(b2, t_36, t_37);
not(t_38, u);
not(t_39, g1);
and(c2, t_38, t_39);
not(t_40, s);
not(t_41, g1);
and(d2, t_40, t_41);
not(t_42, r);
not(t_43, h1);
or(e2, t_42, t_43);
not(t_44, q);
not(t_45, i1);
and(f2, t_44, t_45);
not(t_46, o);
not(t_47, i1);
and(g2, t_46, t_47);
not(t_48, n);
not(t_49, j1);
or(h2, t_48, t_49);
not(t_50, m);
not(t_51, k1);
and(i2, t_50, t_51);
not(t_52, k);
not(t_53, k1);
and(j2, t_52, t_53);
not(t_54, j);
not(t_55, l1);
or(k2, t_54, t_55);
not(t_56, i);
not(t_57, m1);
and(l2, t_56, t_57);
not(t_58, g);
not(t_59, m1);
and(m2, t_58, t_59);
not(t_60, f);
not(t_61, n1);
or(n2, t_60, t_61);
not(t_62, e);
not(t_63, o1);
and(o2, t_62, t_63);
not(t_64, c);
not(t_65, o1);
and(p2, t_64, t_65);
not(t_66, b);
not(t_67, p1);
or(q2, t_66, t_67);
and(r2, q2, n2, k2, h2, e2, b2, y1, v1, s1);
not(s2, r2);
not(t2, r2);
not(t_68, s1);
not(t_69, s2);
and(t_70, s2, t_68);
and(t_71, t_69, s1);
or(u2, t_70, t_71);
not(t_72, f0);
not(t_73, t2);
or(v2, t_72, t_73);
not(t_74, v1);
not(t_75, s2);
and(t_76, s2, t_74);
and(t_77, t_75, v1);
or(w2, t_76, t_77);
not(t_78, b0);
not(t_79, t2);
or(x2, t_78, t_79);
not(t_80, y1);
not(t_81, s2);
and(t_82, s2, t_80);
and(t_83, t_81, y1);
or(y2, t_82, t_83);
not(t_84, x);
not(t_85, t2);
or(z2, t_84, t_85);
not(t_86, b2);
not(t_87, s2);
and(t_88, s2, t_86);
and(t_89, t_87, b2);
or(a3, t_88, t_89);
not(t_90, t);
not(t_91, t2);
or(b3, t_90, t_91);
not(t_92, e2);
not(t_93, s2);
and(t_94, s2, t_92);
and(t_95, t_93, e2);
or(c3, t_94, t_95);
not(t_96, p);
not(t_97, t2);
or(d3, t_96, t_97);
not(t_98, h2);
not(t_99, s2);
and(t_100, s2, t_98);
and(t_101, t_99, h2);
or(e3, t_100, t_101);
not(t_102, l);
not(t_103, t2);
or(f3, t_102, t_103);
not(t_104, k2);
not(t_105, s2);
and(t_106, s2, t_104);
and(t_107, t_105, k2);
or(g3, t_106, t_107);
not(t_108, h);
not(t_109, t2);
or(h3, t_108, t_109);
not(t_110, n2);
not(t_111, s2);
and(t_112, s2, t_110);
and(t_113, t_111, n2);
or(i3, t_112, t_113);
not(t_114, d);
not(t_115, t2);
or(j3, t_114, t_115);
not(t_116, q2);
not(t_117, s2);
and(t_118, s2, t_116);
and(t_119, t_117, q2);
or(k3, t_118, t_119);
not(t_120, t2);
not(t_121, a);
or(l3, t_120, t_121);
not(t_122, q1);
not(t_123, u2);
or(m3, t_122, t_123);
not(t_124, r1);
not(t_125, u2);
or(n3, t_124, t_125);
not(t_126, t1);
not(t_127, w2);
or(o3, t_126, t_127);
not(t_128, u1);
not(t_129, w2);
or(p3, t_128, t_129);
not(t_130, w1);
not(t_131, y2);
or(q3, t_130, t_131);
not(t_132, x1);
not(t_133, y2);
or(r3, t_132, t_133);
not(t_134, z1);
not(t_135, a3);
or(s3, t_134, t_135);
not(t_136, a2);
not(t_137, a3);
or(t3, t_136, t_137);
not(t_138, c2);
not(t_139, c3);
or(u3, t_138, t_139);
not(t_140, d2);
not(t_141, c3);
or(v3, t_140, t_141);
not(t_142, f2);
not(t_143, e3);
or(w3, t_142, t_143);
not(t_144, g2);
not(t_145, e3);
or(x3, t_144, t_145);
not(t_146, i2);
not(t_147, g3);
or(y3, t_146, t_147);
not(t_148, j2);
not(t_149, g3);
or(z3, t_148, t_149);
not(t_150, l2);
not(t_151, i3);
or(a4, t_150, t_151);
not(t_152, m2);
not(t_153, i3);
or(b4, t_152, t_153);
not(t_154, o2);
not(t_155, k3);
or(c4, t_154, t_155);
not(t_156, p2);
not(t_157, k3);
or(d4, t_156, t_157);
not(e4, m3);
and(f4, d4, b4, z3, x3, v3, t3, r3, p3, n3);
not(g4, o3);
not(h4, q3);
not(i4, s3);
not(j4, u3);
not(k4, w3);
not(l4, y3);
not(m4, a4);
not(n4, c4);
not(o4, f4);
not(p4, f4);
not(t_158, i0);
not(t_159, p4);
or(q4, t_158, t_159);
not(t_160, n3);
not(t_161, o4);
and(t_162, o4, t_160);
and(t_163, t_161, n3);
or(r4, t_162, t_163);
not(t_164, e0);
not(t_165, p4);
or(s4, t_164, t_165);
not(t_166, p3);
not(t_167, o4);
and(t_168, o4, t_166);
and(t_169, t_167, p3);
or(t4, t_168, t_169);
not(t_170, a0);
not(t_171, p4);
or(u4, t_170, t_171);
not(t_172, r3);
not(t_173, o4);
and(t_174, o4, t_172);
and(t_175, t_173, r3);
or(v4, t_174, t_175);
not(t_176, w);
not(t_177, p4);
or(w4, t_176, t_177);
not(t_178, t3);
not(t_179, o4);
and(t_180, o4, t_178);
and(t_181, t_179, t3);
or(x4, t_180, t_181);
not(t_182, s);
not(t_183, p4);
or(y4, t_182, t_183);
not(t_184, v3);
not(t_185, o4);
and(t_186, o4, t_184);
and(t_187, t_185, v3);
or(z4, t_186, t_187);
not(t_188, o);
not(t_189, p4);
or(a5, t_188, t_189);
not(t_190, x3);
not(t_191, o4);
and(t_192, o4, t_190);
and(t_193, t_191, x3);
or(b5, t_192, t_193);
not(t_194, k);
not(t_195, p4);
or(c5, t_194, t_195);
not(t_196, z3);
not(t_197, o4);
and(t_198, o4, t_196);
and(t_199, t_197, z3);
or(d5, t_198, t_199);
not(t_200, g);
not(t_201, p4);
or(e5, t_200, t_201);
not(t_202, b4);
not(t_203, o4);
and(t_204, o4, t_202);
and(t_205, t_203, b4);
or(f5, t_204, t_205);
not(t_206, p4);
not(t_207, c);
or(g5, t_206, t_207);
not(t_208, d4);
not(t_209, o4);
and(t_210, o4, t_208);
and(t_211, t_209, d4);
or(h5, t_210, t_211);
not(t_212, e4);
not(t_213, r4);
or(i5, t_212, t_213);
not(t_214, g4);
not(t_215, t4);
or(j5, t_214, t_215);
not(t_216, h4);
not(t_217, v4);
or(k5, t_216, t_217);
not(t_218, i4);
not(t_219, x4);
or(l5, t_218, t_219);
not(t_220, j4);
not(t_221, z4);
or(m5, t_220, t_221);
not(t_222, k4);
not(t_223, b5);
or(n5, t_222, t_223);
not(t_224, l4);
not(t_225, d5);
or(o5, t_224, t_225);
not(t_226, m4);
not(t_227, f5);
or(p5, t_226, t_227);
not(t_228, n4);
not(t_229, h5);
or(q5, t_228, t_229);
and(r5, q5, p5, o5, n5, m5, l5, k5, j5, i5);
not(s5, r5);
not(t_230, j0);
not(t_231, s5);
or(t5, t_230, t_231);
not(t_232, g0);
not(t_233, s5);
or(u5, t_232, t_233);
not(t_234, c0);
not(t_235, s5);
or(v5, t_234, t_235);
not(t_236, y);
not(t_237, s5);
or(w5, t_236, t_237);
not(t_238, u);
not(t_239, s5);
or(x5, t_238, t_239);
not(t_240, q);
not(t_241, s5);
or(y5, t_240, t_241);
not(t_242, m);
not(t_243, s5);
or(z5, t_242, t_243);
not(t_244, i);
not(t_245, s5);
or(a6, t_244, t_245);
not(t_246, s5);
not(t_247, e);
or(b6, t_246, t_247);
not(t_248, h0);
not(t_249, t5);
not(t_250, q4);
not(t_251, v2);
or(c6, t_248, t_249, t_250, t_251);
not(t_252, d0);
not(t_253, u5);
not(t_254, s4);
not(t_255, x2);
or(d6, t_252, t_253, t_254, t_255);
not(t_256, z);
not(t_257, v5);
not(t_258, u4);
not(t_259, z2);
or(e6, t_256, t_257, t_258, t_259);
not(t_260, v);
not(t_261, w5);
not(t_262, w4);
not(t_263, b3);
or(f6, t_260, t_261, t_262, t_263);
not(t_264, r);
not(t_265, x5);
not(t_266, y4);
not(t_267, d3);
or(g6, t_264, t_265, t_266, t_267);
not(t_268, n);
not(t_269, y5);
not(t_270, a5);
not(t_271, f3);
or(h6, t_268, t_269, t_270, t_271);
not(t_272, j);
not(t_273, z5);
not(t_274, c5);
not(t_275, h3);
or(i6, t_272, t_273, t_274, t_275);
not(t_276, f);
not(t_277, a6);
not(t_278, e5);
not(t_279, j3);
or(j6, t_276, t_277, t_278, t_279);
not(t_280, b6);
not(t_281, g5);
not(t_282, l3);
not(t_283, b);
or(k6, t_280, t_281, t_282, t_283);
and(l6, j6, i6, h6, g6, f6, e6, d6, c6);
not(m6, d6);
not(n6, e6);
not(o6, f6);
not(p6, h6);
not(q6, k6);
not(t_284, m6);
not(t_285, e6);
not(t_286, h6);
not(t_287, i6);
or(r6, t_284, t_285, t_286, t_287);
not(t_288, g6);
not(t_289, o6);
not(t_290, h6);
not(t_291, i6);
or(s6, t_288, t_289, t_290, t_291);
not(t_292, n6);
not(t_293, h6);
not(t_294, g6);
or(t6, t_292, t_293, t_294);
not(t_295, p6);
not(t_296, i6);
or(u6, t_295, t_296);
endmodule
module top;
	parameter in_width = 36,
		patterns = 5000,
		step = 1;
	reg [1:in_width] in_mem[1:patterns];
	integer index;

	wire i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,
		i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,
		i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,
		i30,i31,i32,i33,i34,i35;

	assign {i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,
		i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,
		i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,
		i30,i31,i32,i33,i34,i35} = 
		$getpattern(in_mem[index]);

	initial $monitor($time,,o0,o1,o2,o3,o4,o5,o6);
	initial
		begin
			$readmemb("patt.mem", in_mem);
			for(index = 1; index <= patterns; index = index + 1)
				#step;
		end

	foobar cct(o0,o1,o2,o3,o4,o5,o6,i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,
		i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,
		i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,
		i30,i31,i32,i33,i34,i35);
endmodule
