// C5315
module foobar(w5, x5, y5, z5, a6, b6, c6, d6, e6, f6, g6, h6, i6, j6, k6, l6, m6, n6, o6, p6, q6, r6, s6, t6, u6, v6, w6, x6, y6, z6, a7, b7, c7, d7, e7, f7, g7, h7, i7, j7, k7, l7, m7, n7, o7, p7, q7, r7, s7, t7, u7, v7, w7, x7, y7, z7, a8, b8, c8, d8, e8, f8, g8, h8, i8, j8, k8, l8, m8, n8, o8, p8, q8, r8, s8, t8, u8, v8, w8, x8, y8, z8, a9, b9, c9, d9, e9, f9, g9, h9, i9, j9, k9, l9, m9, n9, o9, p9, q9, r9, s9, t9, u9, v9, w9, x9, y9, z9, a10, b10, c10, d10, e10, f10, g10, h10, i10, j10, k10, l10, m10, n10, o10, a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2, b2, c2, d2, e2, f2, g2, h2, i2, j2, k2, l2, m2, n2, o2, p2, q2, r2, s2, t2, u2, v2, w2, x2, y2, z2, a3, b3, c3, d3, e3, f3, g3, h3, i3, j3, k3, l3, m3, n3, o3, p3, q3, r3, s3, t3, u3, v3, w3, x3, y3, z3, a4, b4, c4, d4, e4, f4, g4, h4, i4, j4, k4, l4, m4, n4, o4, p4, q4, r4, s4, t4, u4, v4, w4, x4, y4, z4, a5, b5, c5, d5, e5, f5, g5, h5, i5, j5, k5, l5, m5, n5, o5, p5, q5, r5, s5, t5, u5, v5);
input a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2, b2, c2, d2, e2, f2, g2, h2, i2, j2, k2, l2, m2, n2, o2, p2, q2, r2, s2, t2, u2, v2, w2, x2, y2, z2, a3, b3, c3, d3, e3, f3, g3, h3, i3, j3, k3, l3, m3, n3, o3, p3, q3, r3, s3, t3, u3, v3, w3, x3, y3, z3, a4, b4, c4, d4, e4, f4, g4, h4, i4, j4, k4, l4, m4, n4, o4, p4, q4, r4, s4, t4, u4, v4, w4, x4, y4, z4, a5, b5, c5, d5, e5, f5, g5, h5, i5, j5, k5, l5, m5, n5, o5, p5, q5, r5, s5, t5, u5, v5;
output w5, x5, y5, z5, a6, b6, c6, d6, e6, f6, g6, h6, i6, j6, k6, l6, m6, n6, o6, p6, q6, r6, s6, t6, u6, v6, w6, x6, y6, z6, a7, b7, c7, d7, e7, f7, g7, h7, i7, j7, k7, l7, m7, n7, o7, p7, q7, r7, s7, t7, u7, v7, w7, x7, y7, z7, a8, b8, c8, d8, e8, f8, g8, h8, i8, j8, k8, l8, m8, n8, o8, p8, q8, r8, s8, t8, u8, v8, w8, x8, y8, z8, a9, b9, c9, d9, e9, f9, g9, h9, i9, j9, k9, l9, m9, n9, o9, p9, q9, r9, s9, t9, u9, v9, w9, x9, y9, z9, a10, b10, c10, d10, e10, f10, g10, h10, i10, j10, k10, l10, m10, n10, o10;
not(z5, u4);
not(a6, w3);
not(b6, a4);
and(c6, w4, z4);
not(d6, v4);
not(e6, u4);
not(f6, u4);
not(g6, u3);
not(h6, y3);
and(i6, n1, o1);
not(j6, u2);
not(k6, w4);
not(l6, z4);
not(m6, y4);
not(n6, f21);
and(o6, k1, p15);
not(p6, c32);
not(q6, g17);
not(w6, u6);
not(t_0, m1);
not(t_1, b21);
or(x6, t_0, t_1);
not(y6, b21);
not(e7, d7);
not(f7, i49);
not(g7, j49);
not(h7, k49);
not(i7, l49);
and(j7, p43, v30);
and(k7, q43, v30);
and(l7, o43, v30);
and(m7, r43, v30);
and(n7, l62, m60, s52);
and(o7, z60, o61, e61);
and(p7, z64, u65);
and(q7, u68, z67);
and(r7, w68, k68);
and(s7, r64, v65);
or(v7, k75, v71);
or(w7, b77, t73);
or(x7, e75, u71);
or(y7, f77, u73);
not(z7, q77);
not(a8, n83);
not(b8, o83);
not(c8, o86);
or(d8, s31, g39, t83, t77);
not(e8, g85);
not(f8, a85);
not(g8, f85);
or(h8, t31, h39, s83, s77);
not(i8, e85);
not(j8, b85);
not(k8, c85);
not(l8, d85);
and(o8, u81, y82, x82, b83, q82, p84, w86, e88, f88);
and(p8, g74, j81, d82, f82, g82, i84, p86, y87, z87);
and(q8, e87, x30);
and(r8, f87, y30);
or(s8, a32, a39, q85, r85);
or(t8, e32, q38, s85, v85);
or(u8, f32, r38, t85, w85);
or(v8, p31, u38, u85, u83);
or(w8, z31, z38, m85, j85);
or(x8, d32, p38, n85, k85);
or(y8, g32, s38, o85, l85);
or(z8, o31, t38, p85, r83);
and(a9, p88, w30);
and(b9, s88, x30);
and(c9, t88, x30);
and(d9, w88, x30);
and(e9, q88, z30);
and(f9, r88, y30);
and(g9, u88, y30);
and(h9, v88, y30);
and(i9, a31, d90);
or(j9, m89, a90);
not(k9, e90);
not(l9, f90);
not(m9, x88);
not(n9, h87);
and(o9, h17, j89, u2);
not(p9, g90);
not(q9, h90);
not(r9, y88);
not(s9, g87);
or(t9, c31, h38, m90, k90);
or(u9, d31, i38, o90, q90);
or(v9, w31, y38, p90, r90);
or(w9, f31, k38, d89, e89);
or(x9, x31, m38, o87, p87);
or(y9, v31, x38, n90, l90);
or(z9, e31, j38, c89, b89);
or(a10, y31, l38, n87, m87);
and(b10, c90, w30);
and(c10, i91, w30);
and(d10, w91, w30);
and(e10, x91, w30);
and(f10, b90, z30);
and(g10, j91, z30);
and(h10, v91, z30);
and(i10, y91, z30);
or(j10, i21, y37, p97, i90);
or(k10, k21, a38, q97, j90);
or(l10, q31, f39, h98, i98);
or(m10, r31, e39, g98, f98);
not(n10, p98);
not(o10, q98);
buf(r14, u5);
buf(s14, u5);
buf(t14, u5);
buf(u14, u5);
buf(v14, u5);
buf(w14, t5);
buf(x14, t5);
buf(y14, t5);
buf(z14, t5);
buf(a15, t5);
buf(b15, s5);
buf(c15, s5);
buf(d15, r5);
buf(e15, r5);
buf(f15, q5);
buf(g15, q5);
buf(h15, p5);
buf(i15, p5);
not(j15, o5);
not(k15, n5);
not(l15, m5);
not(m15, l5);
not(n15, k5);
not(o15, j5);
not(p15, i5);
not(q15, h5);
not(r15, g5);
buf(s15, g5);
not(t15, f5);
buf(u15, e5);
buf(v15, e5);
buf(w15, d5);
buf(x15, d5);
buf(y15, c5);
buf(z15, c5);
buf(a16, b5);
buf(b16, b5);
not(c16, a5);
buf(u6, v4);
buf(e16, t4);
buf(f16, t4);
buf(g16, s4);
buf(h16, s4);
buf(i16, r4);
buf(j16, r4);
buf(k16, q4);
buf(l16, q4);
buf(m16, p4);
buf(n16, p4);
buf(o16, o4);
buf(p16, o4);
buf(q16, n4);
buf(r16, n4);
buf(s16, m4);
buf(t16, m4);
buf(u16, l4);
buf(v16, l4);
buf(w16, k4);
buf(x16, k4);
buf(y16, j4);
buf(z16, j4);
buf(a17, i4);
buf(b17, i4);
buf(c17, h4);
buf(d17, h4);
buf(e17, g4);
buf(f17, g4);
and(g17, f4, x4);
and(h17, f4, y4, x4, w4);
buf(i17, e4);
buf(j17, e4);
buf(k17, b4);
buf(l17, z3);
buf(m17, z3);
buf(n17, z3);
buf(o17, x3);
buf(p17, x3);
buf(q17, x3);
buf(r17, x3);
buf(s17, x3);
buf(t17, v3);
buf(u17, v3);
buf(v17, v3);
buf(w17, v3);
buf(x17, v3);
buf(y17, t3);
buf(z17, t3);
buf(a18, s3);
buf(b18, s3);
buf(c18, q3);
buf(d18, q3);
buf(e18, q3);
buf(f18, q3);
not(g18, q3);
buf(h18, o3);
buf(i18, o3);
buf(j18, o3);
buf(k18, o3);
buf(l18, o3);
buf(m18, m3);
buf(n18, m3);
buf(o18, m3);
buf(p18, m3);
buf(q18, m3);
buf(r18, k3);
buf(s18, k3);
buf(t18, k3);
buf(v6, j3);
buf(v18, i3);
buf(w18, i3);
buf(x18, i3);
buf(y18, g3);
buf(z18, e3);
buf(a19, e3);
buf(b19, e3);
buf(c19, e3);
buf(d19, e3);
buf(e19, c3);
buf(f19, c3);
buf(g19, c3);
buf(h19, c3);
buf(i19, c3);
buf(j19, a3);
buf(k19, a3);
buf(l19, a3);
buf(m19, a3);
buf(n19, a3);
buf(o19, y2);
buf(p19, y2);
buf(q19, y2);
buf(r19, y2);
buf(s19, y2);
buf(t19, x2);
buf(u19, x2);
buf(v19, w2);
buf(w19, w2);
buf(x19, v2);
buf(y19, v2);
buf(z19, t2);
buf(a20, t2);
buf(b20, r2);
buf(c20, r2);
buf(d20, r2);
buf(e20, r2);
buf(f20, r2);
buf(g20, p2);
buf(h20, p2);
buf(i20, p2);
buf(j20, p2);
buf(k20, p2);
buf(l20, n2);
buf(m20, n2);
buf(n20, n2);
buf(o20, n2);
buf(p20, n2);
buf(q20, l2);
buf(r20, l2);
buf(s20, l2);
buf(t20, l2);
buf(u20, l2);
buf(v20, j2);
buf(s6, n1);
buf(r6, l1);
buf(y20, l1);
and(z20, j1, v5);
buf(a21, u);
and(b21, k, l);
and(c21, l, k);
buf(d21, b);
buf(t6, a);
not(t_2, a);
not(t_3, d4);
or(f21, t_2, t_3);
not(g21, r14);
not(h21, s14);
and(i21, y14, t14);
not(j21, t14);
and(k21, z14, u14);
not(l21, u14);
not(m21, v14);
not(n21, w14);
not(o21, x14);
not(p21, y14);
not(q21, z14);
not(r21, a15);
not(s21, b15);
not(t21, c15);
not(u21, d15);
not(v21, e15);
not(w21, f15);
not(x21, g15);
not(y21, h15);
not(z21, i15);
and(a22, o15, t20);
and(b22, o15, o20);
and(c22, o15, j20);
and(d22, o15, f20);
and(e22, o15, r19);
and(f22, o15, m19);
and(g22, o15, g19);
and(h22, o15, c19);
and(i22, o15, e18);
and(j22, o15, v17);
and(k22, o15, r17);
not(l22, r15);
not(m22, s15);
not(n22, u15);
not(o22, v15);
not(p22, w15);
not(q22, x15);
not(r22, y15);
not(s22, z15);
not(t22, a16);
not(u22, b16);
and(v22, y19, t4, o17);
and(w22, l15, t4, q17);
not(x22, e16);
not(y22, f16);
and(z22, l15, s4, w17);
and(a23, y19, s4, u17);
not(b23, g16);
not(c23, h16);
or(d23, r4, a20);
and(e23, y19, r4);
or(f23, r4, o15);
and(g23, l15, r4);
not(h23, i16);
not(i23, j16);
and(j23, l15, q4, f18);
and(k23, y19, q4, d18);
not(l23, k16);
not(m23, l16);
and(n23, y19, p4, h18);
and(o23, x19, p4, j18);
not(p23, m16);
not(q23, n16);
and(r23, x19, o4, q18);
and(s23, y19, o4, o18);
not(t23, o16);
not(u23, p16);
and(v23, x19, n4, l20);
and(w23, l15, n4, n20);
not(x23, q16);
not(y23, r16);
and(z23, x19, m4, s20);
and(a24, l15, m4, u20);
not(b24, s16);
not(c24, t16);
not(d24, u16);
not(e24, v16);
and(f24, x19, k4, b20);
and(g24, l15, k4, e20);
not(h24, w16);
not(i24, x16);
and(j24, x19, j4, i20);
and(k24, l15, j4, k20);
not(l24, y16);
not(m24, z16);
and(n24, l15, i4, h19);
and(o24, x19, i4, f19);
not(p24, a17);
not(q24, b17);
and(r24, x19, h4, j19);
and(s24, l15, h4, l19);
not(t24, c17);
not(u24, d17);
and(v24, l15, g4, s19);
and(w24, x19, g4, q19);
not(x24, e17);
not(y24, f17);
and(z24, x19, e4, z18);
and(a25, l15, e4, b19);
not(b25, i17);
not(c25, j17);
and(d25, c4, b18);
not(e25, k17);
and(f25, a4, b18);
and(g25, y19, l17);
not(h25, l17);
and(i25, y19, m17);
not(j25, m17);
not(k25, n17);
and(l25, y3, b18);
not(m25, o17);
and(n25, a20, p17);
not(o25, p17);
not(p25, q17);
not(q25, r17);
not(r25, s17);
and(s25, w3, b18);
and(t25, a20, t17);
not(u25, t17);
not(v25, u17);
not(w25, v17);
not(x25, w17);
not(y25, x17);
and(z25, u3, b18);
not(a26, y17);
not(b26, z17);
not(c26, a18);
not(d26, b18);
and(e26, r3, a18);
and(f26, a20, c18);
not(g26, c18);
not(h26, d18);
not(i26, e18);
not(j26, f18);
buf(k26, g18);
buf(l26, g18);
and(m26, p3, a18);
not(n26, h18);
and(o26, a20, i18);
not(p26, i18);
not(q26, j18);
and(r26, z19, k18);
not(s26, k18);
not(t26, l18);
and(u26, n3, a18);
not(v26, m18);
and(w26, a20, n18);
not(x26, n18);
not(y26, o18);
and(z26, z19, p18);
not(a27, p18);
not(b27, q18);
and(c27, l3, a18);
and(d27, y19, r18);
not(e27, r18);
not(f27, s18);
and(g27, x19, t18);
not(h27, t18);
buf(d7, v6);
and(j27, j3, a18);
not(k27, v18);
and(l27, a20, w18);
not(m27, w18);
and(n27, z19, x18);
not(o27, x18);
and(p27, h3, z17);
not(q27, y18);
and(r27, f3, z17);
not(s27, z18);
and(t27, z19, a19);
not(u27, a19);
not(v27, b19);
not(w27, c19);
not(x27, d19);
and(y27, d3, z17);
and(z27, z19, e19);
not(a28, e19);
not(b28, f19);
not(c28, g19);
not(d28, h19);
not(e28, i19);
and(f28, b3, z17);
not(g28, j19);
and(h28, z19, k19);
not(i28, k19);
not(j28, l19);
not(k28, m19);
not(l28, n19);
and(m28, z2, z17);
not(n28, o19);
and(o28, z19, p19);
not(p28, p19);
not(q28, q19);
not(r28, r19);
not(s28, s19);
and(t28, z19, r20);
and(u28, z19, m20);
and(v28, z19, h20);
and(w28, z19, c20);
and(x28, s2, y17);
not(y28, b20);
not(z28, c20);
not(a29, d20);
not(b29, e20);
not(c29, f20);
and(d29, q2, y17);
not(e29, g20);
not(f29, h20);
not(g29, i20);
not(h29, j20);
not(i29, k20);
and(j29, o2, y17);
not(k29, l20);
not(l29, m20);
not(m29, n20);
not(n29, o20);
not(o29, p20);
and(p29, m2, y17);
not(q29, q20);
not(r29, r20);
not(s29, s20);
not(t29, t20);
not(u29, u20);
and(v29, k2, y17);
buf(w29, v20);
buf(x29, v20);
buf(y29, v20);
buf(z29, v20);
buf(a30, v20);
and(b30, c2, a16, y15);
and(c30, c2, w15, u15);
and(d30, a2, a16, y15);
and(e30, a2, w15, u15);
and(f30, y1, x15, v15);
and(g30, y1, b16, z15);
and(h30, x1, b16, z15);
and(i30, x1, x15, v15);
and(j30, w1, b16, z15);
and(k30, w1, x15, v15);
and(l30, v1, x15, v15);
and(m30, v1, b16, z15);
and(n30, u1, b16, z15);
and(o30, u1, x15, v15);
and(p30, t1, w15, u15);
and(q30, t1, a16, y15);
and(r30, r1, a16, y15);
and(s30, r1, w15, u15);
and(t30, p1, w15, u15);
and(u30, p1, a16, y15);
buf(v30, s6);
buf(w30, r6);
buf(x30, r6);
buf(y30, y20);
buf(z30, y20);
not(a31, z20);
and(b31, b1, j15, n5);
and(c31, o0, d15, b15);
and(d31, o0, f15, h15);
and(e31, n0, d15, b15);
and(f31, n0, f15, h15);
and(g31, l0, v14);
and(h31, l0, v14);
and(i31, k0, v14);
and(j31, k0, v14);
and(k31, i0, r15);
and(l31, i0, r15);
and(m31, g0, r15);
and(n31, f0, r15);
and(o31, y, e15, c15);
and(p31, y, g15, i15);
and(q31, w, g15, i15);
and(r31, w, e15, c15);
and(s31, v, g15, i15);
and(t31, v, e15, c15);
not(u31, a21);
and(v31, r, d15, b15);
and(w31, r, f15, h15);
and(x31, o, f15, h15);
and(y31, o, d15, b15);
and(z31, n, d15, b15);
and(a32, n, f15, h15);
not(b32, b21);
and(c32, q15, k);
and(d32, f, e15, c15);
and(e32, f, g15, i15);
and(f32, e, g15, i15);
and(g32, e, e15, c15);
not(h32, d21);
buf(i32, t6);
and(j32, n15, t29);
and(k32, n15, n29);
and(l32, n15, h29);
and(m32, n15, c29);
and(n32, n15, r28);
and(o32, n15, k28);
and(p32, n15, c28);
and(q32, n15, w27);
and(r32, n15, i26);
and(s32, n15, w25);
and(t32, n15, q25);
and(u32, s15, b32);
and(v32, s15, b32);
and(w32, s15, b32);
and(x32, s15, b32);
and(y32, m22, b32);
and(z32, m22, b32);
and(a33, m22, b32);
and(b33, m22, b32);
and(c33, t4, w19, m25);
and(d33, t4, m15, p25);
and(e33, s4, m15, x25);
and(f33, s4, w19, v25);
not(g33, e23);
not(h33, g23);
and(i33, q4, m15, j26);
and(j33, q4, w19, h26);
and(k33, p4, w19, n26);
and(l33, p4, v19, q26);
and(m33, o4, v19, b27);
and(n33, o4, w19, y26);
and(o33, n4, v19, k29);
and(p33, n4, m15, m29);
and(q33, m4, v19, s29);
and(r33, m4, m15, u29);
and(s33, y19, l4, z29);
and(t33, y19, l4, x29);
and(u33, k4, v19, y28);
and(v33, k4, m15, b29);
and(w33, j4, v19, g29);
and(x33, j4, m15, i29);
and(y33, i4, m15, d28);
and(z33, i4, v19, b28);
and(a34, h4, v19, g28);
and(b34, h4, m15, j28);
and(c34, g4, m15, s28);
and(d34, g4, v19, q28);
and(e34, e4, v19, s27);
and(f34, e4, m15, v27);
and(g34, b4, d26);
not(t_4, k25);
not(t_5, k17);
or(h34, t_4, t_5);
and(i34, z3, d26);
not(t_6, e25);
not(t_7, n17);
or(j34, t_6, t_7);
and(k34, x3, d26);
not(t_8, y25);
not(t_9, s17);
or(l34, t_8, t_9);
and(m34, v3, d26);
not(t_10, r25);
not(t_11, x17);
or(n34, t_10, t_11);
or(o34, z25, d26);
and(p34, q3, c26);
not(q34, k26);
not(r34, l26);
and(s34, o3, c26);
not(t_12, v26);
not(t_13, l18);
or(t34, t_12, t_13);
not(t_14, t26);
not(t_15, m18);
or(u34, t_14, t_15);
and(v34, m3, c26);
not(t_16, k27);
not(t_17, s18);
or(w34, t_16, t_17);
and(x34, k3, c26);
not(t_18, f27);
not(t_19, v18);
or(y34, t_18, t_19);
and(z34, i3, c26);
and(a35, g3, b26);
not(t_20, x27);
not(t_21, y18);
or(b35, t_20, t_21);
and(c35, e3, b26);
not(t_22, q27);
not(t_23, d19);
or(d35, t_22, t_23);
and(e35, c3, b26);
not(t_24, l28);
not(t_25, i19);
or(f35, t_24, t_25);
and(g35, a3, b26);
not(t_26, e28);
not(t_27, n19);
or(h35, t_26, t_27);
not(t_28, a29);
not(t_29, o19);
or(i35, t_28, t_29);
and(j35, y2, b26);
and(k35, t19, o27);
and(l35, t19, a27);
and(m35, t19, s26);
and(n35, t19, p28);
and(o35, t19, i28);
and(p35, t19, a28);
and(q35, t19, u27);
and(r35, t19, r29);
and(s35, t19, l29);
and(t35, t19, f29);
and(u35, t19, z28);
and(v35, u19, g26);
and(w35, u19, o25);
and(x35, u19, u25);
and(y35, u19, m27);
and(z35, u19, p26);
and(a36, u19, x26);
and(b36, v19, h27);
and(c36, w19, h25);
and(d36, w19, j25);
and(e36, w19, e27);
and(f36, a20, w29);
and(g36, a20, y29);
and(h36, r2, a26);
not(t_30, n28);
not(t_31, d20);
or(i36, t_30, t_31);
not(t_32, o29);
not(t_33, g20);
or(j36, t_32, t_33);
and(k36, p2, a26);
and(l36, n2, a26);
not(t_34, e29);
not(t_35, p20);
or(m36, t_34, t_35);
not(t_36, q29);
not(t_37, a30);
or(n36, t_36, t_37);
and(o36, l2, a26);
not(p36, w29);
not(q36, x29);
not(r36, y29);
not(s36, z29);
not(t36, a30);
and(u36, j2, a26);
and(v36, i2, q22, v15);
and(w36, i2, u22, z15);
and(x36, h2, q22, v15);
and(y36, h2, u22, z15);
and(z36, g2, q22, v15);
and(a37, g2, u22, z15);
and(b37, f2, q22, v15);
and(c37, f2, u22, z15);
and(d37, e2, q22, v15);
and(e37, e2, u22, z15);
and(f37, d2, t22, y15);
and(g37, d2, p22, u15);
and(h37, b2, p22, u15);
and(i37, b2, t22, y15);
and(j37, z1, p22, u15);
and(k37, z1, t22, y15);
and(l37, s1, p22, u15);
and(m37, s1, t22, y15);
and(n37, q1, t22, y15);
and(o37, q1, p22, u15);
and(p37, h1, p21, t14);
and(q37, g1, p21, t14);
and(r37, f1, p21, t14);
and(s37, e1, q21, u14);
and(t37, d1, q21, u14);
and(u37, c1, q21, u14);
and(v37, b1, n21, r14);
and(w37, a1, o21, s14);
and(x37, z0, n21, r14);
and(y37, y0, p21, t14);
and(z37, x0, p21, t14);
and(a38, w0, q21, u14);
and(b38, v0, q21, u14);
and(c38, u0, n21, r14);
and(d38, t0, o21, s14);
and(e38, s0, o21, s14);
and(f38, r0, o21, s14);
and(g38, q0, n21, r14);
and(h38, p0, u21, b15);
and(i38, p0, w21, h15);
and(j38, m0, u21, b15);
and(k38, m0, w21, h15);
and(l38, j0, u21, b15);
and(m38, j0, w21, h15);
and(n38, h0, l22);
and(o38, f0, l22);
and(p38, a0, v21, c15);
and(q38, a0, x21, i15);
and(r38, z, x21, i15);
and(s38, z, v21, c15);
and(t38, x, v21, c15);
and(u38, x, x21, i15);
and(v38, t, o21, s14);
and(w38, s, n21, r14);
and(x38, q, u21, b15);
and(y38, q, w21, h15);
and(z38, p, u21, b15);
and(a39, p, w21, h15);
and(b39, m, l22);
and(c39, m, l22);
not(d39, b32);
and(e39, d, v21, c15);
and(f39, d, x21, i15);
and(g39, c, x21, i15);
and(h39, c, v21, c15);
or(i39, t4, w35, n25);
or(j39, c33, v22);
or(k39, t4, t32, k22);
or(l39, d33, w22);
or(m39, e33, z22);
or(n39, s4, s32, j22);
or(o39, f33, a23);
or(p39, s4, x35, t25);
and(q39, g33, d23);
and(r39, h33, f23);
and(s39, r4, o34);
and(t39, o34, r4);
or(u39, i33, j23);
or(v39, q4, r32, i22);
or(w39, j33, k23);
or(x39, q4, v35, f26);
or(y39, p4, z35, o26);
or(z39, k33, n23);
or(a40, p4, m35, r26);
or(b40, l33, o23);
or(c40, m33, r23);
or(d40, o4, l35, z26);
or(e40, n33, s23);
or(f40, o4, a36, w26);
or(g40, n4, s35, u28);
or(h40, o33, v23);
or(i40, n4, k32, b22);
or(j40, p33, w23);
or(k40, q33, z23);
or(l40, m4, r35, t28);
or(m40, r33, a24);
or(n40, m4, j32, a22);
and(o40, l4, w19, s36);
and(p40, l4, w19, q36);
or(q40, k4, u35, w28);
or(r40, u33, f24);
or(s40, k4, m32, d22);
or(t40, v33, g24);
or(u40, w33, j24);
or(v40, j4, t35, v28);
or(w40, x33, k24);
or(x40, j4, l32, c22);
or(y40, y33, n24);
or(z40, i4, p32, g22);
or(a41, z33, o24);
or(b41, i4, p35, z27);
or(c41, h4, o35, h28);
or(d41, a34, r24);
or(e41, h4, o32, f22);
or(f41, b34, s24);
or(g41, c34, v24);
or(h41, g4, n32, e22);
or(i41, d34, w24);
or(j41, g4, n35, o28);
or(k41, e4, q35, t27);
or(l41, e34, z24);
or(m41, e4, q32, h22);
or(n41, f34, a25);
or(o41, d25, g34);
not(t_38, j34);
not(t_39, h34);
or(p41, t_38, t_39);
or(q41, f25, i34);
or(r41, c36, g25);
or(s41, d36, i25);
or(t41, l25, k34);
not(t_40, n34);
not(t_41, l34);
or(u41, t_40, t_41);
or(v41, s25, m34);
buf(w41, o34);
buf(x41, o34);
buf(y41, o34);
or(z41, e26, p34);
or(a42, m26, s34);
not(t_42, u34);
not(t_43, t34);
or(b42, t_42, t_43);
or(c42, u26, v34);
or(d42, c27, x34);
or(e42, e36, d27);
not(t_44, y34);
not(t_45, w34);
or(f42, t_44, t_45);
or(g42, b36, g27);
or(h42, j27, z34);
or(i42, y35, l27);
or(j42, k35, n27);
or(k42, p27, a35);
not(t_46, d35);
not(t_47, b35);
or(l42, t_46, t_47);
or(m42, r27, c35);
or(n42, y27, e35);
not(t_48, h35);
not(t_49, f35);
or(o42, t_48, t_49);
or(p42, f28, g35);
or(q42, m28, j35);
not(t_50, i36);
not(t_51, i35);
or(r42, t_50, t_51);
and(s42, u19, p36);
and(t42, u19, r36);
or(u42, x28, h36);
or(v42, d29, k36);
not(t_52, m36);
not(t_53, j36);
or(w42, t_52, t_53);
or(x42, j29, l36);
or(y42, p29, o36);
not(t_54, t36);
not(t_55, q20);
or(z42, t_54, t_55);
or(a43, v29, u36);
or(b43, k31, b39);
or(c43, l31, c39);
or(d43, m31, n38);
or(e43, n31, o38);
and(f43, e0, m22, d39);
and(g43, d0, s15, d39);
and(h43, c0, s15, d39);
and(i43, b0, m22, d39);
and(j43, j, m22, d39);
and(k43, i, s15, d39);
and(l43, h, m22, d39);
and(m43, g, s15, d39);
and(n43, r39, p21, j21);
or(o43, u32, y32, m43, i43);
or(p43, v32, b33, k43, l43);
or(q43, w32, a33, g43, j43);
or(r43, x32, z32, h43, f43);
not(s43, j39);
not(t43, l39);
and(u43, t4, t41);
and(v43, t41, t4);
not(w43, m39);
not(x43, o39);
and(y43, v41, s4);
and(z43, s4, v41);
not(a44, q39);
not(b44, r39);
not(t_56, h23);
not(t_57, x41);
or(c44, t_56, t_57);
not(t_58, i23);
not(t_59, w41);
or(d44, t_58, t_59);
not(e44, u39);
not(f44, w39);
and(g44, q4, z41);
and(h44, z41, q4);
not(i44, z39);
not(j44, b40);
not(t_60, p4);
not(t_61, a42);
and(k44, t_60, t_61);
and(l44, p4, a42);
and(m44, p4, a42);
not(t_62, p4);
not(t_63, a42);
and(n44, t_62, t_63);
not(o44, c40);
not(p44, e40);
and(q44, c42, o4);
and(r44, o4, c42);
not(s44, h40);
not(t44, j40);
and(u44, x42, n4);
and(v44, n4, x42);
not(w44, k40);
not(x44, m40);
and(y44, m4, y42);
and(z44, y42, m4);
or(a45, l4, t42, g36);
or(b45, o40, s33);
or(c45, l4, s42, f36);
or(d45, p40, t33);
and(e45, a43, l4);
and(f45, l4, a43);
not(g45, r40);
not(h45, t40);
and(i45, k4, u42);
and(j45, u42, k4);
not(k45, u40);
not(l45, w40);
and(m45, j4, v42);
not(t_64, j4);
not(t_65, v42);
and(n45, t_64, t_65);
not(t_66, j4);
not(t_67, v42);
and(o45, t_66, t_67);
and(p45, j4, v42);
not(q45, y40);
not(r45, a41);
and(s45, n42, i4);
and(t45, i4, n42);
not(u45, d41);
not(v45, f41);
and(w45, h4, p42);
and(x45, p42, h4);
not(y45, g41);
not(z45, i41);
and(a46, q42, g4);
and(b46, g4, q42);
not(c46, l41);
not(d46, n41);
not(t_68, e4);
not(t_69, m42);
and(e46, t_68, t_69);
and(f46, e4, m42);
and(g46, m42, e4);
not(h46, o41);
not(i46, p41);
not(j46, q41);
buf(k46, q41);
buf(l46, q41);
not(m46, q41);
buf(n46, q41);
not(o46, r41);
not(p46, s41);
buf(q46, t41);
buf(r46, t41);
buf(s46, t41);
not(t46, u41);
buf(u46, v41);
buf(v46, v41);
buf(w46, v41);
not(x46, w41);
not(y46, x41);
not(z46, y41);
buf(a47, z41);
buf(b47, z41);
buf(c47, z41);
and(d47, u41, p41, l26);
buf(e47, a42);
buf(f47, a42);
buf(g47, a42);
not(h47, b42);
buf(i47, c42);
buf(j47, c42);
buf(k47, c42);
not(l47, d42);
buf(m47, d42);
not(n47, d42);
buf(o47, d42);
buf(p47, d42);
not(q47, e42);
not(r47, f42);
not(s47, g42);
not(t47, h42);
not(u47, h42);
buf(v47, h42);
buf(w47, h42);
not(x47, i42);
not(y47, j42);
buf(z47, j42);
not(a48, k42);
not(b48, l42);
buf(c48, m42);
buf(d48, m42);
buf(e48, m42);
buf(f48, n42);
buf(g48, n42);
buf(h48, n42);
not(i48, o42);
buf(j48, p42);
buf(k48, p42);
buf(l48, p42);
buf(m48, q42);
buf(n48, q42);
buf(o48, q42);
buf(p48, r42);
buf(q48, r42);
buf(r48, u42);
buf(s48, u42);
buf(t48, u42);
buf(u48, v42);
buf(v48, v42);
buf(w48, v42);
not(x48, w42);
buf(y48, x42);
buf(z48, x42);
buf(a49, x42);
buf(b49, y42);
buf(c49, y42);
buf(d49, y42);
not(t_70, n36);
not(t_71, z42);
or(e49, t_70, t_71);
buf(f49, a43);
buf(g49, a43);
buf(h49, a43);
and(i49, d43, c21);
and(j49, c43, c21);
and(k49, b43, c21);
and(l49, e43, c21);
and(m49, s47, n21, g21);
and(n49, z47, n21, g21);
and(o49, o46, p21, j21);
and(p49, z47, j15, k15);
and(q49, s43, i39);
and(r49, t43, k39);
not(t_72, x22);
not(t_73, r46);
or(s49, t_72, t_73);
not(t_74, y22);
not(t_75, q46);
or(t49, t_74, t_75);
and(u49, w43, n39);
and(v49, x43, p39);
not(t_76, b23);
not(t_77, w46);
or(w49, t_76, t_77);
not(t_78, c23);
not(t_79, v46);
or(x49, t_78, t_79);
not(t_80, y46);
not(t_81, i16);
or(y49, t_80, t_81);
not(t_82, x46);
not(t_83, j16);
or(z49, t_82, t_83);
and(a50, e44, v39);
and(b50, f44, x39);
not(t_84, l23);
not(t_85, c47);
or(c50, t_84, t_85);
not(t_86, m23);
not(t_87, b47);
or(d50, t_86, t_87);
and(e50, i44, y39);
and(f50, j44, a40);
not(t_88, p23);
not(t_89, f47);
or(g50, t_88, t_89);
not(h50, k44);
buf(i50, l44);
not(t_90, q23);
not(t_91, g47);
or(j50, t_90, t_91);
buf(k50, m44);
not(l50, n44);
and(m50, o44, d40);
and(n50, p44, f40);
not(t_92, t23);
not(t_93, j47);
or(o50, t_92, t_93);
and(p50, l47, t47, q44);
and(q50, l47, q44);
and(r50, l47, q44);
not(t_94, u23);
not(t_95, k47);
or(s50, t_94, t_95);
and(t50, n47, r44);
and(u50, n47, u47, r44);
and(v50, n47, r44);
and(w50, s44, g40);
and(x50, t44, i40);
not(t_96, x23);
not(t_97, z48);
or(y50, t_96, t_97);
not(t_98, y23);
not(t_99, a49);
or(z50, t_98, t_99);
and(a51, w44, l40);
and(b51, x44, n40);
not(t_100, b24);
not(t_101, c49);
or(c51, t_100, t_101);
not(t_102, c24);
not(t_103, d49);
or(d51, t_102, t_103);
not(e51, b45);
not(f51, d45);
not(t_104, d24);
not(t_105, g49);
or(g51, t_104, t_105);
not(t_106, e24);
not(t_107, h49);
or(h51, t_106, t_107);
and(i51, g45, q40);
and(j51, h45, s40);
not(t_108, h24);
not(t_109, t48);
or(k51, t_108, t_109);
not(t_110, i24);
not(t_111, s48);
or(l51, t_110, t_111);
and(m51, k45, v40);
and(n51, l45, x40);
not(t_112, l24);
not(t_113, w48);
or(o51, t_112, t_113);
buf(p51, m45);
not(q51, n45);
not(t_114, m24);
not(t_115, v48);
or(r51, t_114, t_115);
not(s51, o45);
buf(t51, p45);
and(u51, q45, z40);
and(v51, r45, b41);
not(t_116, p24);
not(t_117, h48);
or(w51, t_116, t_117);
not(t_118, q24);
not(t_119, g48);
or(x51, t_118, t_119);
and(y51, u45, c41);
and(z51, v45, e41);
not(t_120, t24);
not(t_121, l48);
or(a52, t_120, t_121);
not(t_122, u24);
not(t_123, k48);
or(b52, t_122, t_123);
and(c52, y45, h41);
and(d52, z45, j41);
not(t_124, x24);
not(t_125, o48);
or(e52, t_124, t_125);
not(t_126, y24);
not(t_127, n48);
or(f52, t_126, t_127);
and(g52, c46, k41);
and(h52, d46, m41);
not(t_128, b25);
not(t_129, e48);
or(i52, t_128, t_129);
not(j52, e46);
buf(k52, f46);
not(t_130, c25);
not(t_131, d48);
or(l52, t_130, t_131);
not(t_132, h46);
not(t_133, n46);
or(m52, t_132, t_133);
buf(n52, j46);
buf(o52, l46);
buf(p52, m46);
buf(q52, m46);
not(r52, n46);
not(s52, p46);
not(t52, p46);
not(u52, q46);
not(v52, r46);
not(w52, s46);
not(x52, u46);
not(y52, v46);
not(z52, w46);
not(t_134, z46);
not(t_135, a47);
or(a53, t_134, t_135);
not(b53, a47);
not(c53, b47);
not(d53, c47);
and(e53, t46, i46, k26);
and(f53, p41, t46, q34);
and(g53, i46, u41, r34);
not(h53, e47);
not(i53, f47);
not(j53, g47);
not(t_136, r47);
not(t_137, b42);
or(k53, t_136, t_137);
not(l53, i47);
not(m53, j47);
not(n53, k47);
buf(o53, l47);
buf(p53, l47);
and(q53, t47, m47);
buf(r53, n47);
buf(s53, n47);
and(t53, u47, o47);
not(u53, p47);
not(t_138, x47);
not(t_139, q47);
or(v53, t_138, t_139);
not(w53, q47);
not(t_140, h47);
not(t_141, f42);
or(x53, t_140, t_141);
not(y53, s47);
buf(z53, t47);
buf(a54, t47);
buf(b54, u47);
buf(c54, u47);
not(d54, v47);
not(e54, w47);
not(t_142, a48);
not(t_143, f49);
or(f54, t_142, t_143);
and(g54, o42, l42, p48);
and(h54, i48, b48, q48);
not(i54, c48);
not(j54, d48);
not(k54, e48);
not(l54, f48);
not(m54, g48);
not(n54, h48);
not(o54, j48);
not(p54, k48);
not(q54, l48);
not(r54, m48);
not(s54, n48);
not(t54, o48);
not(u54, p48);
not(v54, q48);
not(w54, r48);
not(x54, s48);
not(y54, t48);
not(z54, u48);
not(a55, v48);
not(b55, w48);
not(t_144, x48);
not(t_145, e49);
or(c55, t_144, t_145);
not(d55, y48);
not(e55, z48);
not(f55, a49);
not(g55, b49);
not(h55, c49);
not(i55, d49);
not(j55, e49);
not(k55, f49);
not(l55, g49);
not(m55, h49);
and(n55, u, j46);
and(o55, a50, n21, g21);
and(p55, f50, n21, g21);
and(q55, m50, n21, g21);
and(r55, j51, o21, h21);
and(s55, n51, o21, h21);
and(t55, x50, o21, h21);
and(u55, b51, o21, h21);
and(v55, r49, p21, j21);
and(w55, u49, p21, j21);
and(x55, h52, q21, l21);
and(y55, u51, q21, l21);
and(z55, z51, q21, l21);
and(a56, c52, q21, l21);
not(b56, q49);
not(c56, r49);
not(t_146, v52);
not(t_147, e16);
or(d56, t_146, t_147);
not(t_148, u52);
not(t_149, f16);
or(e56, t_148, t_149);
not(f56, u49);
not(g56, v49);
not(t_150, z52);
not(t_151, g16);
or(h56, t_150, t_151);
not(t_152, y52);
not(t_153, h16);
or(i56, t_152, t_153);
not(t_154, a44);
not(t_155, b50);
or(j56, t_154, t_155);
not(t_156, y49);
not(t_157, c44);
or(k56, t_156, t_157);
not(t_158, d44);
not(t_159, z49);
or(l56, t_158, t_159);
not(m56, a50);
not(n56, b50);
not(t_160, d53);
not(t_161, k16);
or(o56, t_160, t_161);
not(t_162, c53);
not(t_163, l16);
or(p56, t_162, t_163);
not(q56, e50);
not(r56, f50);
not(t_164, i53);
not(t_165, m16);
or(s56, t_164, t_165);
not(t56, i50);
not(t_166, j53);
not(t_167, n16);
or(u56, t_166, t_167);
not(v56, k50);
not(w56, m50);
not(x56, n50);
not(t_168, m53);
not(t_169, o16);
or(y56, t_168, t_169);
not(t_170, n53);
not(t_171, p16);
or(z56, t_170, t_171);
not(a57, w50);
not(b57, x50);
not(t_172, e55);
not(t_173, q16);
or(c57, t_172, t_173);
not(t_174, f55);
not(t_175, r16);
or(d57, t_174, t_175);
not(e57, a51);
not(f57, b51);
not(t_176, h55);
not(t_177, s16);
or(g57, t_176, t_177);
not(t_178, i55);
not(t_179, t16);
or(h57, t_178, t_179);
and(i57, e51, a45);
and(j57, f51, c45);
not(t_180, l55);
not(t_181, u16);
or(k57, t_180, t_181);
not(t_182, m55);
not(t_183, v16);
or(l57, t_182, t_183);
not(m57, i51);
not(n57, j51);
not(t_184, y54);
not(t_185, w16);
or(o57, t_184, t_185);
not(t_186, x54);
not(t_187, x16);
or(p57, t_186, t_187);
not(q57, m51);
not(r57, n51);
not(t_188, b55);
not(t_189, y16);
or(s57, t_188, t_189);
not(t57, p51);
not(t_190, a55);
not(t_191, z16);
or(u57, t_190, t_191);
not(v57, t51);
not(w57, u51);
not(x57, v51);
not(t_192, n54);
not(t_193, a17);
or(y57, t_192, t_193);
not(t_194, m54);
not(t_195, b17);
or(z57, t_194, t_195);
not(a58, y51);
not(b58, z51);
not(t_196, q54);
not(t_197, c17);
or(c58, t_196, t_197);
not(t_198, p54);
not(t_199, d17);
or(d58, t_198, t_199);
not(e58, c52);
not(f58, d52);
not(t_200, t54);
not(t_201, e17);
or(g58, t_200, t_201);
not(t_202, s54);
not(t_203, f17);
or(h58, t_202, t_203);
not(i58, g52);
not(j58, h52);
not(t_204, k54);
not(t_205, i17);
or(k58, t_204, t_205);
not(l58, k52);
not(t_206, j54);
not(t_207, j17);
or(m58, t_206, t_207);
not(t_208, r52);
not(t_209, o41);
or(n58, t_208, t_209);
not(o58, n52);
or(p58, n55, k46);
not(q58, o52);
not(r58, p52);
not(s58, q52);
not(t58, t52);
not(t_210, x52);
not(t_211, s46);
or(u58, t_210, t_211);
not(t_212, w52);
not(t_213, u46);
or(v58, t_212, t_213);
not(t_214, b53);
not(t_215, y41);
or(w58, t_214, t_215);
not(t_216, f53);
not(t_217, e53);
and(x58, t_216, t_217);
not(t_218, g53);
not(t_219, d47);
and(y58, t_218, t_219);
not(t_220, l53);
not(t_221, e47);
or(z58, t_220, t_221);
not(t_222, x53);
not(t_223, k53);
or(a59, t_222, t_223);
not(t_224, h53);
not(t_225, i47);
or(b59, t_224, t_225);
not(c59, o53);
not(d59, p53);
not(e59, r53);
not(f59, s53);
not(t_226, d54);
not(t_227, p47);
or(g59, t_226, t_227);
not(h59, z53);
not(i59, a54);
not(j59, b54);
not(k59, c54);
not(t_228, u53);
not(t_229, v47);
or(l59, t_228, t_229);
and(m59, e54, w47);
not(t_230, w53);
not(t_231, i42);
or(n59, t_230, t_231);
not(t_232, k55);
not(t_233, k42);
or(o59, t_232, t_233);
and(p59, l42, i48, v54);
not(t_234, l54);
not(t_235, c48);
or(q59, t_234, t_235);
not(t_236, i54);
not(t_237, f48);
or(r59, t_236, t_237);
and(s59, b48, o42, u54);
not(t_238, r54);
not(t_239, j48);
or(t59, t_238, t_239);
not(t_240, o54);
not(t_241, m48);
or(u59, t_240, t_241);
not(t_242, z54);
not(t_243, r48);
or(v59, t_242, t_243);
not(t_244, w54);
not(t_245, u48);
or(w59, t_244, t_245);
not(t_246, j55);
not(t_247, w42);
or(x59, t_246, t_247);
not(t_248, g55);
not(t_249, y48);
or(y59, t_248, t_249);
not(t_250, d55);
not(t_251, b49);
or(z59, t_250, t_251);
not(t_252, u31);
not(t_253, n52);
or(a60, t_252, t_253);
and(b60, i57, o21, h21);
not(t_254, g56);
not(t_255, q49);
or(c60, t_254, t_255);
not(t_256, d56);
not(t_257, s49);
or(d60, t_256, t_257);
not(t_258, t49);
not(t_259, e56);
or(e60, t_258, t_259);
not(t_260, b56);
not(t_261, v49);
or(f60, t_260, t_261);
not(t_262, w49);
not(t_263, h56);
or(g60, t_262, t_263);
and(h60, l56, y43);
not(t_264, i56);
not(t_265, x49);
or(i60, t_264, t_265);
and(j60, k56, z43);
and(k60, k56, z43);
not(t_266, n56);
not(t_267, q39);
or(l60, t_266, t_267);
and(m60, c56, f56, b44, m56);
buf(n60, k56);
buf(o60, k56);
buf(p60, l56);
not(t_268, o56);
not(t_269, c50);
or(q60, t_268, t_269);
not(t_270, d50);
not(t_271, p56);
or(r60, t_270, t_271);
not(t_272, x56);
not(t_273, e50);
or(s60, t_272, t_273);
not(t_274, s56);
not(t_275, g50);
or(t60, t_274, t_275);
not(t_276, j50);
not(t_277, u56);
or(u60, t_276, t_277);
not(t_278, q56);
not(t_279, n50);
or(v60, t_278, t_279);
not(t_280, o50);
not(t_281, y56);
or(w60, t_280, t_281);
not(t_282, z56);
not(t_283, s50);
or(x60, t_282, t_283);
not(t_284, q57);
not(t_285, w50);
or(y60, t_284, t_285);
and(z60, n57, r57, b57, f57);
not(t_286, y50);
not(t_287, c57);
or(a61, t_286, t_287);
not(t_288, d57);
not(t_289, z50);
or(b61, t_288, t_289);
not(t_290, g57);
not(t_291, c51);
or(c61, t_290, t_291);
not(t_292, d51);
not(t_293, h57);
or(d61, t_292, t_293);
not(e61, j57);
buf(f61, j57);
not(t_294, g51);
not(t_295, k57);
or(g61, t_294, t_295);
not(t_296, l57);
not(t_297, h51);
or(h61, t_296, t_297);
not(t_298, f58);
not(t_299, i51);
or(i61, t_298, t_299);
not(t_300, o57);
not(t_301, k51);
or(j61, t_300, t_301);
not(t_302, l51);
not(t_303, p57);
or(k61, t_302, t_303);
not(t_304, a57);
not(t_305, m51);
or(l61, t_304, t_305);
not(t_306, o51);
not(t_307, s57);
or(m61, t_306, t_307);
not(t_308, u57);
not(t_309, r51);
or(n61, t_308, t_309);
and(o61, j58, w57, b58, e58);
not(t_310, a58);
not(t_311, v51);
or(p61, t_310, t_311);
not(t_312, w51);
not(t_313, y57);
or(q61, t_312, t_313);
not(t_314, z57);
not(t_315, x51);
or(r61, t_314, t_315);
not(t_316, x57);
not(t_317, y51);
or(s61, t_316, t_317);
not(t_318, c58);
not(t_319, a52);
or(t61, t_318, t_319);
not(t_320, b52);
not(t_321, d58);
or(u61, t_320, t_321);
not(t_322, m57);
not(t_323, d52);
or(v61, t_322, t_323);
not(t_324, e52);
not(t_325, g58);
or(w61, t_324, t_325);
not(t_326, h58);
not(t_327, f52);
or(x61, t_326, t_327);
not(y61, i58);
not(t_328, k58);
not(t_329, i52);
or(z61, t_328, t_329);
not(t_330, l52);
not(t_331, m58);
or(a62, t_330, t_331);
not(t_332, n58);
not(t_333, m52);
or(b62, t_332, t_333);
not(c62, p58);
not(t_334, u58);
not(t_335, v58);
or(d62, t_334, t_335);
not(t_336, a53);
not(t_337, w58);
or(e62, t_336, t_337);
not(t_338, y58);
not(t_339, x58);
or(f62, t_338, t_339);
not(t_340, b59);
not(t_341, z58);
or(g62, t_340, t_341);
not(h62, a59);
not(t_342, l59);
not(t_343, g59);
or(i62, t_342, t_343);
not(t_344, n59);
not(t_345, v53);
or(j62, t_344, t_345);
or(k62, m59, e54);
and(l62, r56, w56, y53, y47);
not(t_346, o59);
not(t_347, f54);
or(m62, t_346, t_347);
not(t_348, s59);
not(t_349, g54);
and(n62, t_348, t_349);
not(t_350, p59);
not(t_351, h54);
and(o62, t_350, t_351);
not(t_352, r59);
not(t_353, q59);
or(p62, t_352, t_353);
not(t_354, u59);
not(t_355, t59);
or(q62, t_354, t_355);
not(t_356, w59);
not(t_357, v59);
or(r62, t_356, t_357);
not(t_358, c55);
not(t_359, x59);
or(s62, t_358, t_359);
not(t_360, z59);
not(t_361, y59);
or(t62, t_360, t_361);
not(t_362, o58);
not(t_363, a21);
or(u62, t_362, t_363);
not(t_364, f60);
not(t_365, c60);
or(v62, t_364, t_365);
buf(w62, d60);
buf(x62, d60);
and(y62, i60, u43, k56);
and(z62, i60, u43, k56);
and(a63, i60, q60, u43, k56);
and(b63, i60, u43);
and(c63, i60, u43);
and(d63, g60, v43, l56);
and(e63, g60, r60, v43, l56);
and(f63, v43, g60);
buf(g63, e60);
buf(h63, g60);
and(i63, l56, r60, y43);
buf(j63, i60);
buf(k63, i60);
and(l63, k56, q60, z43);
not(t_366, j56);
not(t_367, l60);
or(m63, t_366, t_367);
not(n63, n60);
not(o63, o60);
and(p63, q60, s39);
not(q63, p60);
and(r63, r60, t39);
buf(s63, q60);
buf(t63, q60);
buf(u63, r60);
not(t_368, v60);
not(t_369, s60);
or(v63, t_368, t_369);
buf(w63, t60);
and(x63, t60, x60);
buf(y63, t60);
and(z63, x60, l44, n47);
and(a64, x60, u47, l44, n47);
and(b64, x60, l44, n47);
and(c64, x60, l44);
and(d64, u60, w60);
not(e64, u60);
and(f64, w60, t47, m44, l47);
and(g64, m44, w60, l47);
and(h64, w60, m44, l47);
and(i64, w60, m44);
and(j64, w60, m44);
buf(k64, w60);
buf(l64, w60);
buf(m64, x60);
buf(n64, x60);
not(t_370, y60);
not(t_371, l61);
or(o64, t_370, t_371);
buf(p64, a61);
buf(q64, a61);
and(r64, d61, m61, a61, g61);
and(s64, m61, a61, d61);
and(t64, m61, a61);
and(u64, d61, g61, u44);
and(v64, d61, u44);
and(w64, d61, u44);
and(x64, n61, b61);
buf(y64, b61);
and(z64, n61, b61, c61, h61);
and(a65, n61, b61, c61);
buf(b65, b61);
and(c65, c61, v44);
and(d65, c61, h61, v44);
and(e65, c61, v44);
not(t_372, e57);
not(t_373, f61);
or(f65, t_372, t_373);
buf(g65, c61);
buf(h65, c61);
and(i65, h61, y44);
buf(j65, d61);
buf(k65, d61);
and(l65, g61, z44);
not(m65, f61);
buf(n65, g61);
buf(o65, g61);
buf(p65, h61);
buf(q65, h61);
not(t_374, i61);
not(t_375, v61);
or(r65, t_374, t_375);
buf(s65, j61);
buf(t65, j61);
and(u65, z61, r61, t61, x61, j61);
and(v65, w61, a62, u61, k61, q61);
buf(w65, k61);
not(x65, m61);
and(y65, a61, g61, m45, d61);
and(z65, m45, a61, d61);
and(a66, a61, m45, d61);
and(b66, a61, m45);
and(c66, a61, m45);
buf(d66, n61);
buf(e66, n61);
and(f66, b61, p45, c61);
and(g66, b61, h61, p45, c61);
and(h66, b61, p45, c61);
and(i66, b61, p45);
not(t_376, s61);
not(t_377, p61);
or(j66, t_376, t_377);
and(k66, u61, s45, w61);
and(l66, u61, k61, s45, w61);
and(m66, s45, u61);
buf(n66, q61);
buf(o66, r61);
and(p66, z61, t61, x61, r61);
and(q66, z61, t61, r61);
buf(r66, r61);
and(s66, z61, r61);
and(t66, t61, t45, x61);
and(u66, t61, t45, x61);
and(v66, t61, j61, t45, x61);
and(w66, t61, t45);
and(x66, t61, t45);
buf(y66, t61);
buf(z66, t61);
and(a67, x61, w45);
and(b67, x61, w45);
and(c67, x61, j61, w45);
buf(d67, u61);
and(e67, w61, x45);
and(f67, w61, k61, x45);
buf(g67, w61);
and(h67, k61, a46);
buf(i67, x61);
buf(j67, x61);
and(k67, j61, b46);
buf(l67, z61);
buf(m67, z61);
and(n67, r61, t61, f46, x61);
and(o67, r61, t61, j61, f46, x61);
and(p67, r61, t61, f46, x61);
and(q67, r61, t61, f46);
and(r67, r61, f46);
and(s67, r61, t61, f46);
buf(t67, a62);
and(u67, q61, u61, g46, w61);
and(v67, q61, u61, k61, g46, w61);
and(w67, q61, g46);
and(x67, q61, u61, g46);
not(y67, b62);
and(z67, l56, j46, g60, r60, e60);
and(a68, e60, g60, k46, l56);
and(b68, e60, g60, r60, k46, l56);
and(c68, e60, k46);
and(d68, e60, g60, k46);
and(e68, d60, i60, l46, k56);
and(f68, d60, i60, q60, l46, k56);
and(g68, d60, i60, l46, k56);
and(h68, d60, i60, l46);
and(i68, d60, l46);
and(j68, d60, i60, l46);
and(k68, m46, d60, i60, k56, q60);
and(l68, m46, i60, k56, d60);
and(m68, m46, d60);
and(n68, m46, i60, d60);
not(o68, d62);
buf(p68, e62);
buf(q68, e62);
not(t_378, h62);
not(t_379, f62);
or(r68, t_378, t_379);
not(s68, f62);
not(t68, g62);
and(u68, l47, u60, w60, t47);
and(v68, u60, w60, l47);
and(w68, t60, x60, n47, u47);
and(x68, t60, x60, n47);
not(y68, i62);
not(z68, j62);
buf(a69, m62);
buf(b69, m62);
not(t_380, n62);
not(t_381, o62);
or(c69, t_380, t_381);
not(d69, p62);
not(e69, q62);
not(f69, r62);
not(g69, s62);
not(h69, t62);
not(t_382, i1);
not(t_383, k62);
or(i69, t_382, t_383);
and(j69, u, j46, g60, e60, l56);
and(k69, u, j46, e60);
not(t_384, u62);
not(t_385, a60);
or(l69, t_384, t_385);
and(m69, u, j46, g60, e60);
and(n69, b, a62, u61, q61, w61);
and(o69, b, a62);
and(p69, b, a62, q61);
and(q69, b, a62, u61, q61);
and(r69, l69, y14, j21);
not(s69, v62);
not(t69, w62);
not(u69, x62);
or(v69, i68, u43);
or(w69, k69, c68, v43);
not(x69, g63);
not(y69, h63);
or(z69, m69, d68, f63, y43);
not(a70, j63);
not(b70, k63);
not(t_386, z43);
not(t_387, b63);
not(t_388, j68);
and(c70, t_386, t_387, t_388);
or(d70, n68, h68, c63, z43);
buf(e70, m63);
buf(f70, m63);
not(t_389, s39);
not(t_390, j60);
not(t_391, y62);
not(t_392, g68);
and(g70, t_389, t_390, t_391, t_392);
or(h70, l68, e68, z62, k60, s39);
or(i70, j69, a68, d63, h60, t39);
not(j70, s63);
not(k70, t63);
or(l70, f68, a63, l63, p63, g44);
not(m70, u63);
or(n70, b68, e63, i63, r63, h44);
not(t_393, z68);
not(t_394, v63);
or(o70, t_393, t_394);
not(p70, v63);
not(q70, w63);
not(r70, y63);
not(t_395, v56);
not(t_396, k64);
or(s70, t_395, t_396);
not(t_397, l50);
not(t_398, l64);
or(t70, t_397, t_398);
not(u70, k64);
not(v70, l64);
not(t_399, q44);
not(t_400, j64);
and(w70, t_399, t_400);
or(x70, d64, i64, q44);
not(y70, m64);
not(z70, n64);
or(a71, c64, r44);
not(b71, o64);
not(c71, p64);
not(d71, q64);
not(t_401, u44);
not(t_402, c66);
and(e71, t_401, t_402);
or(f71, t64, b66, u44);
not(g71, y64);
not(h71, b65);
or(i71, i66, v44);
not(t_403, m65);
not(t_404, a51);
or(j71, t_403, t_404);
not(k71, g65);
not(l71, h65);
not(t_405, y44);
not(t_406, c65);
not(t_407, h66);
and(m71, t_405, t_406, t_407);
or(n71, a65, f66, e65, y44);
not(o71, j65);
not(p71, k65);
not(t_408, z44);
not(t_409, w64);
not(t_410, z65);
and(q71, t_408, t_409, t_410);
or(r71, s64, a66, v64, z44);
not(s71, n65);
not(t71, o65);
or(u71, y65, u64, l65, e45);
or(v71, g66, d65, i65, f45);
not(w71, p65);
not(x71, q65);
buf(y71, r65);
buf(z71, r65);
not(a72, s65);
not(b72, t65);
not(c72, u65);
or(d72, o67, v66, c67, k67, i45);
not(e72, w65);
or(f72, v67, l66, f67, h67, j45);
not(t_411, t57);
not(t_412, p64);
or(g72, t_411, t_412);
not(t_413, q51);
not(t_414, q64);
or(h72, t_413, t_414);
not(i72, d66);
not(j72, e66);
not(k72, j66);
or(l72, p69, w67, s45);
not(m72, n66);
not(n72, o66);
not(o72, r66);
or(p72, r67, t45);
not(q72, y66);
not(r72, z66);
not(t_415, w45);
not(t_416, w66);
not(t_417, s67);
and(s72, t_415, t_416, t_417);
or(t72, q66, q67, x66, w45);
not(u72, d67);
or(v72, q69, x67, m66, x45);
not(w72, g67);
or(x72, n69, u67, k66, e67, a46);
not(y72, i67);
not(z72, j67);
not(t_418, b46);
not(t_419, a67);
not(t_420, t66);
not(t_421, p67);
and(a73, t_418, t_419, t_420, t_421);
or(b73, p66, n67, u66, b67, b46);
not(c73, l67);
not(d73, m67);
not(e73, t67);
or(f73, o69, g46);
and(g73, b62, d62, q68);
and(h73, y67, o68, p68);
not(t_422, c62);
not(t_423, g63);
or(i73, t_422, t_423);
not(j73, k68);
not(k73, p68);
not(l73, q68);
not(t_424, y68);
not(t_425, g62);
or(m73, t_424, t_425);
not(t_426, s68);
not(t_427, a59);
or(n73, t_426, t_427);
not(t_428, m47);
not(t_429, r50);
not(t_430, g64);
and(o73, t_428, t_429, t_430);
or(p73, v68, h64, q50, m47);
not(t_431, o47);
not(t_432, t50);
not(t_433, b64);
and(q73, t_431, t_432, t_433);
or(r73, x68, z63, v50, o47);
not(t_434, t68);
not(t_435, i62);
or(s73, t_434, t_435);
or(t73, f64, p50, q53, h42);
or(u73, a64, u50, t53, h42);
and(v73, k62, i69);
not(w73, a69);
and(x73, h69, f69, b69);
not(y73, b69);
not(t_436, g69);
not(t_437, c69);
or(z73, t_436, t_437);
not(a74, c69);
not(t_438, e69);
not(t_439, p62);
or(b74, t_438, t_439);
not(t_440, d69);
not(t_441, q62);
or(c74, t_440, t_441);
and(d74, t62, r62, a69);
and(e74, i69, i1);
and(f74, z67, u);
not(g74, l69);
and(h74, v65, b);
not(t_442, h32);
not(t_443, t67);
or(i74, t_442, t_443);
not(j74, v69);
not(t_444, y69);
not(t_445, w69);
or(k74, t_444, t_445);
not(l74, w69);
not(m74, z69);
not(n74, c70);
not(o74, d70);
not(p74, e70);
not(q74, f70);
not(r74, g70);
not(s74, h70);
not(t_446, q63);
not(t_447, z69);
or(t74, t_446, t_447);
not(t_448, m70);
not(t_449, i70);
or(u74, t_448, t_449);
not(v74, i70);
not(w74, l70);
or(x74, f74, n70);
or(y74, x63, a71);
not(t_450, u70);
not(t_451, k50);
or(z74, t_450, t_451);
not(t_452, v70);
not(t_453, n44);
or(a75, t_452, t_453);
not(b75, w70);
not(c75, x70);
not(d75, a71);
and(e75, f72, r64);
not(t_454, o71);
not(t_455, e71);
or(f75, t_454, t_455);
not(g75, e71);
not(t_456, p71);
not(t_457, f71);
or(h75, t_456, t_457);
not(i75, f71);
or(j75, x64, i71);
and(k75, z64, d72);
not(l75, i71);
not(t_458, f65);
not(t_459, j71);
or(m75, t_458, t_459);
not(n75, m71);
not(o75, n71);
not(t_460, t71);
not(t_461, q71);
or(p75, t_460, t_461);
not(q75, q71);
not(t_462, s71);
not(t_463, r71);
or(r75, t_462, t_463);
not(s75, r71);
not(t75, y71);
not(u75, z71);
not(v75, d72);
not(t_464, e72);
not(t_465, x72);
or(w75, t_464, t_465);
or(x75, h74, f72);
not(t_466, c71);
not(t_467, p51);
or(y75, t_466, t_467);
not(t_468, d71);
not(t_469, n45);
or(z75, t_468, t_469);
not(t_470, u72);
not(t_471, l72);
or(a76, t_470, t_471);
not(b76, l72);
not(t_472, m72);
not(t_473, f73);
or(c76, t_472, t_473);
or(d76, s66, p72);
not(e76, p72);
not(f76, s72);
not(g76, t72);
not(t_474, w72);
not(t_475, v72);
or(h76, t_474, t_475);
not(i76, v72);
not(j76, x72);
not(k76, a73);
not(l76, b73);
and(m76, j66, i58, z71);
and(n76, k72, y61, y71);
not(t_476, j52);
not(t_477, t72);
or(o76, t_476, t_477);
not(t_478, l58);
not(t_479, s72);
or(p76, t_478, t_479);
not(q76, f73);
and(r76, o68, b62, l73);
not(t_480, x69);
not(t_481, p58);
or(s76, t_480, t_481);
not(t_482, q58);
not(t_483, c70);
or(t76, t_482, t_483);
or(u76, m68, v69);
and(v76, v62, t52, f70);
and(w76, s69, t58, e70);
and(x76, d62, y67, k73);
not(t_484, r68);
not(t_485, n73);
or(t7, t_484, t_485);
not(t_486, s73);
not(t_487, m73);
or(z76, t_486, t_487);
not(t_488, c59);
not(t_489, w70);
or(a77, t_488, t_489);
and(b77, n70, u68);
not(t_490, d59);
not(t_491, x70);
or(c77, t_490, t_491);
not(d77, o73);
not(e77, p73);
and(f77, w68, l70);
not(g77, q73);
not(h77, r73);
not(t_492, p70);
not(t_493, j62);
or(i77, t_492, t_493);
not(t_494, h59);
not(t_495, p73);
or(j77, t_494, t_495);
not(t_496, i59);
not(t_497, o73);
or(k77, t_496, t_497);
or(l77, e74, v73);
not(t_498, c74);
not(t_499, b74);
or(m77, t_498, t_499);
and(n77, r62, h69, y73);
not(t_500, a74);
not(t_501, s62);
or(o77, t_500, t_501);
and(p77, f69, t62, w73);
or(q77, p37, r69, o49);
not(t_502, e73);
not(t_503, d21);
or(r77, t_502, t_503);
and(s77, q77, v21, t21);
and(t77, q77, x21, z21);
and(u77, l77, o5, k15);
and(v77, q77, p22, n22);
and(w77, q77, t22, r22);
not(x77, j74);
not(t_504, l74);
not(t_505, h63);
or(y77, t_504, t_505);
not(t_506, o74);
not(t_507, u76);
or(z77, t_506, t_507);
not(t_508, m74);
not(t_509, p60);
or(a78, t_508, t_509);
not(t_510, v74);
not(t_511, u63);
or(b78, t_510, t_511);
not(c78, x74);
not(t_512, i77);
not(t_513, o70);
or(d78, t_512, t_513);
not(e78, y74);
not(t_514, h50);
not(t_515, y74);
or(f78, t_514, t_515);
not(t_516, t56);
not(t_517, d75);
or(g78, t_516, t_517);
and(h78, x74, e64);
not(t_518, z74);
not(t_519, s70);
or(i78, t_518, t_519);
not(t_520, a75);
not(t_521, t70);
or(j78, t_520, t_521);
not(k78, d75);
not(t_522, b71);
not(t_523, m75);
or(l78, t_522, t_523);
not(m78, j75);
not(n78, l75);
not(o78, m75);
not(t_524, g75);
not(t_525, j65);
or(p78, t_524, t_525);
not(t_526, i75);
not(t_527, k65);
or(q78, t_526, t_527);
not(t_528, s75);
not(t_529, n65);
or(r78, t_528, t_529);
not(t_530, q75);
not(t_531, o65);
or(s78, t_530, t_531);
and(t78, v75, c72);
not(t_532, j76);
not(t_533, w65);
or(u78, t_532, t_533);
not(v78, x75);
and(w78, x75, x65);
not(t_534, y75);
not(t_535, g72);
or(x78, t_534, t_535);
not(t_536, z75);
not(t_537, h72);
or(y78, t_536, t_537);
not(t_538, s51);
not(t_539, j75);
or(z78, t_538, t_539);
not(t_540, v57);
not(t_541, l75);
or(a79, t_540, t_541);
not(t_542, q76);
not(t_543, n66);
or(b79, t_542, t_543);
not(c79, d76);
not(d79, e76);
not(t_544, b76);
not(t_545, d67);
or(e79, t_544, t_545);
not(t_546, i76);
not(t_547, g67);
or(f79, t_546, t_547);
and(g79, i58, k72, t75);
and(h79, y61, j66, u75);
not(t_548, g76);
not(t_549, e46);
or(i79, t_548, t_549);
not(t_550, f76);
not(t_551, k52);
or(j79, t_550, t_551);
not(t_552, r76);
not(t_553, g73);
and(k79, t_552, t_553);
not(t_554, x76);
not(t_555, h73);
and(l79, t_554, t_555);
not(t_556, s76);
not(t_557, i73);
or(m79, t_556, t_557);
not(t_558, n74);
not(t_559, o52);
or(n79, t_558, t_559);
and(o79, w74, j73);
not(p79, u76);
and(q79, t52, s69, p74);
and(r79, t58, v62, q74);
not(s79, t7);
not(t79, z76);
not(t_560, b75);
not(t_561, o53);
or(u79, t_560, t_561);
not(t_562, c75);
not(t_563, p53);
or(v79, t_562, t_563);
not(t_564, e77);
not(t_565, z53);
or(w79, t_564, t_565);
not(t_566, d77);
not(t_567, a54);
or(x79, t_566, t_567);
not(t_568, n77);
not(t_569, x73);
and(y79, t_568, t_569);
not(t_570, z73);
not(t_571, o77);
or(u7, t_570, t_571);
not(a80, m77);
not(t_572, p77);
not(t_573, d74);
and(b80, t_572, t_573);
not(t_574, r77);
not(t_575, i74);
or(c80, t_574, t_575);
and(d80, m79, y14, j21);
and(e80, c80, z14, l21);
not(t_576, k74);
not(t_577, y77);
or(f80, t_576, t_577);
not(t_578, p79);
not(t_579, d70);
or(g80, t_578, t_579);
not(t_580, t74);
not(t_581, a78);
or(h80, t_580, t_581);
not(t_582, u74);
not(t_583, b78);
or(i80, t_582, t_583);
and(j80, i78, c78);
not(k80, d78);
not(t_584, e78);
not(t_585, k44);
or(l80, t_584, t_585);
not(t_586, k78);
not(t_587, i50);
or(m80, t_586, t_587);
and(n80, u60, c78);
not(o80, j78);
not(t_588, o78);
not(t_589, o64);
or(p80, t_588, t_589);
not(t_590, f75);
not(t_591, p78);
or(q80, t_590, t_591);
not(t_592, h75);
not(t_593, q78);
or(r80, t_592, t_593);
not(t_594, p75);
not(t_595, s78);
or(s80, t_594, t_595);
not(t_596, r75);
not(t_597, r78);
or(t80, t_596, t_597);
not(u80, t78);
not(t_598, w75);
not(t_599, u78);
or(v80, t_598, t_599);
and(w80, x78, v78);
and(x80, m61, v78);
not(y80, y78);
not(t_600, m78);
not(t_601, o45);
or(z80, t_600, t_601);
not(t_602, n78);
not(t_603, t51);
or(a81, t_602, t_603);
not(t_604, a76);
not(t_605, e79);
or(b81, t_604, t_605);
not(t_606, c76);
not(t_607, b79);
or(c81, t_606, t_607);
not(t_608, h76);
not(t_609, f79);
or(d81, t_608, t_609);
not(t_610, h79);
not(t_611, m76);
and(e81, t_610, t_611);
not(t_612, g79);
not(t_613, n76);
and(f81, t_612, t_613);
not(t_614, i79);
not(t_615, o76);
or(g81, t_614, t_615);
not(t_616, j79);
not(t_617, p76);
or(h81, t_616, t_617);
not(t_618, k79);
not(t_619, l79);
or(i81, t_618, t_619);
not(j81, m79);
not(t_620, n79);
not(t_621, t76);
or(k81, t_620, t_621);
not(l81, o79);
not(t_622, r79);
not(t_623, v76);
and(m81, t_622, t_623);
not(t_624, q79);
not(t_625, w76);
and(n81, t_624, t_625);
not(t_626, a77);
not(t_627, u79);
or(o81, t_626, t_627);
not(t_628, c77);
not(t_629, v79);
or(p81, t_628, t_629);
not(t_630, j77);
not(t_631, w79);
or(q81, t_630, t_631);
not(t_632, k77);
not(t_633, x79);
or(r81, t_632, t_633);
not(t_634, b80);
not(t_635, y79);
or(s81, t_634, t_635);
not(t81, u7);
not(u81, c80);
and(v81, i80, w14, g21);
and(w81, v80, x14, h21);
and(x81, h80, y14, j21);
and(y81, f80, y14, j21);
and(z81, d81, z14, l21);
and(a82, b81, z14, l21);
and(b82, c81, z14, l21);
not(t_636, x77);
not(t_637, k81);
or(c82, t_636, t_637);
not(d82, f80);
not(t_638, g80);
not(t_639, z77);
or(e82, t_638, t_639);
not(f82, h80);
not(g82, i80);
and(h82, x74, p81);
and(i82, x74, o80);
and(j82, x74, q81);
not(t_640, l80);
not(t_641, f78);
or(k82, t_640, t_641);
not(t_642, m80);
not(t_643, g78);
or(l82, t_642, t_643);
or(m82, h78, n80);
not(t_644, l78);
not(t_645, p80);
or(n82, t_644, t_645);
not(o82, q80);
not(p82, s80);
not(q82, v80);
and(r82, x75, r80);
and(s82, x75, y80);
and(t82, x75, t80);
or(u82, w78, x80);
not(t_646, z80);
not(t_647, z78);
or(v82, t_646, t_647);
not(t_648, a81);
not(t_649, a79);
or(w82, t_648, t_649);
not(x82, b81);
not(y82, c81);
not(t_650, c79);
not(t_651, g81);
or(z82, t_650, t_651);
not(t_652, d79);
not(t_653, h81);
or(a83, t_652, t_653);
not(b83, d81);
not(t_654, e81);
not(t_655, f81);
or(c83, t_654, t_655);
not(d83, g81);
not(e83, h81);
not(f83, i81);
not(g83, k81);
not(t_656, m81);
not(t_657, n81);
or(h83, t_656, t_657);
not(t_658, t79);
not(t_659, i81);
or(i83, t_658, t_659);
not(j83, o81);
not(k83, r81);
not(l83, s81);
not(t_660, a80);
not(t_661, s81);
or(m83, t_660, t_661);
or(n83, r37, d80, v55);
or(o83, b38, e80, x55);
and(p83, m82, w14, g21);
and(q83, u82, x14, h21);
and(r83, n83, v21, t21);
and(s83, o83, e15, t21);
and(t83, o83, g15, z21);
and(u83, n83, x21, z21);
and(v83, n83, p22, n22);
and(w83, o83, w15, n22);
and(x83, n83, t22, r22);
and(y83, o83, a16, r22);
not(t_662, g83);
not(t_663, j74);
or(z83, t_662, t_663);
not(a84, e82);
not(t_664, s74);
not(t_665, e82);
or(b84, t_664, t_665);
and(c84, k83, c78);
or(d84, i82, j80);
and(e84, j83, c78);
not(t_666, k80);
not(t_667, h83);
or(f84, t_666, t_667);
not(g84, k82);
not(h84, l82);
not(i84, m82);
not(j84, n82);
not(t_668, n75);
not(t_669, w82);
or(k84, t_668, t_669);
not(t_670, o75);
not(t_671, v82);
or(l84, t_670, t_671);
and(m84, p82, v78);
or(n84, s82, w80);
and(o84, o82, v78);
not(p84, u82);
not(q84, v82);
not(r84, w82);
not(t_672, d83);
not(t_673, d76);
or(s84, t_672, t_673);
not(t_674, e83);
not(t_675, e76);
or(t84, t_674, t_675);
not(u84, c83);
not(v84, h83);
not(t_676, f83);
not(t_677, z76);
or(w84, t_676, t_677);
not(t_678, g77);
not(t_679, l82);
or(x84, t_678, t_679);
not(t_680, h77);
not(t_681, k82);
or(y84, t_680, t_681);
not(t_682, l83);
not(t_683, m77);
or(z84, t_682, t_683);
or(a85, q37, x81, n43);
or(b85, s37, z81, a56);
or(c85, t37, a82, z55);
or(d85, u37, b82, y55);
or(e85, w37, w81, r55);
or(f85, z37, y81, w55);
or(g85, w38, v81, o55);
and(h85, d84, w14, g21);
and(i85, n84, x14, h21);
and(j85, g85, u21, s21);
and(k85, a85, v21, t21);
and(l85, f85, v21, t21);
and(m85, e85, d15, s21);
and(n85, b85, e15, t21);
and(o85, c85, e15, t21);
and(p85, d85, e15, t21);
and(q85, e85, f15, y21);
and(r85, g85, w21, y21);
and(s85, b85, g15, z21);
and(t85, c85, g15, z21);
and(u85, d85, g15, z21);
and(v85, a85, x21, z21);
and(w85, f85, x21, z21);
and(x85, f85, p22, n22);
and(y85, a85, p22, n22);
and(z85, g85, q22, o22);
and(a86, b85, w15, n22);
and(b86, c85, w15, n22);
and(c86, d85, w15, n22);
and(d86, e85, x15, o22);
and(e86, f85, t22, r22);
and(f86, a85, t22, r22);
and(g86, g85, u22, s22);
and(h86, b85, a16, r22);
and(i86, c85, a16, r22);
and(j86, d85, a16, r22);
and(k86, e85, b16, s22);
not(t_684, c82);
not(t_685, z83);
or(l86, t_684, t_685);
not(t_686, a84);
not(t_687, h70);
or(m86, t_686, t_687);
or(n86, h82, e84);
or(o86, j82, c84);
not(p86, d84);
not(t_688, v84);
not(t_689, d78);
or(q86, t_688, t_689);
not(t_690, u84);
not(t_691, n82);
or(r86, t_690, t_691);
not(t_692, r84);
not(t_693, m71);
or(s86, t_692, t_693);
not(t_694, q84);
not(t_695, n71);
or(t86, t_694, t_695);
or(u86, r82, o84);
or(v86, t82, m84);
not(w86, n84);
not(t_696, z82);
not(t_697, s84);
or(x86, t_696, t_697);
not(t_698, a83);
not(t_699, t84);
or(y86, t_698, t_699);
not(t_700, j84);
not(t_701, c83);
or(z86, t_700, t_701);
not(t_702, i83);
not(t_703, w84);
or(m8, t_702, t_703);
not(t_704, h84);
not(t_705, q73);
or(b87, t_704, t_705);
not(t_706, g84);
not(t_707, r73);
or(c87, t_706, t_707);
not(t_708, m83);
not(t_709, z84);
or(n8, t_708, t_709);
or(e87, b30, i37, y83, w77);
or(f87, c30, h37, w83, v77);
or(g87, f38, q83, s55);
or(h87, g38, p83, p55);
and(i87, o86, w14, g21);
and(j87, n86, w14, g21);
and(k87, v86, x14, h21);
and(l87, u86, x14, h21);
and(m87, h87, u21, s21);
and(n87, g87, d15, s21);
and(o87, g87, f15, y21);
and(p87, h87, w21, y21);
and(q87, o86, o5, n5);
and(r87, h87, q22, o22);
and(s87, g87, x15, o22);
and(t87, h87, u22, s22);
and(u87, g87, b16, s22);
not(v87, l86);
not(t_710, r74);
not(t_711, l86);
or(w87, t_710, t_711);
not(t_712, b84);
not(t_713, m86);
or(x87, t_712, t_713);
not(y87, n86);
not(z87, o86);
not(t_714, f84);
not(t_715, q86);
or(a88, t_714, t_715);
not(t_716, z86);
not(t_717, r86);
or(b88, t_716, t_717);
not(t_718, k84);
not(t_719, s86);
or(c88, t_718, t_719);
not(t_720, l84);
not(t_721, t86);
or(d88, t_720, t_721);
not(e88, u86);
not(f88, v86);
not(g88, x86);
not(h88, y86);
not(t_722, k76);
not(t_723, y86);
or(i88, t_722, t_723);
not(t_724, l76);
not(t_725, x86);
or(j88, t_724, t_725);
not(k88, m8);
not(t_726, x84);
not(t_727, b87);
or(l88, t_726, t_727);
not(t_728, y84);
not(t_729, c87);
or(m88, t_728, t_729);
not(t_730, o86);
not(t_731, l77);
or(n88, t_730, t_731);
not(o88, n8);
or(p88, h30, y36, k86, g86);
or(q88, i30, x36, d86, z85);
or(r88, p30, g37, c86, v83);
or(s88, q30, f37, j86, x83);
or(t88, r30, m37, i86, e86);
or(u88, s30, l37, b86, x85);
or(v88, t30, o37, a86, y85);
or(w88, u30, n37, h86, f86);
or(x88, c38, h85, q55);
or(y88, v38, i85, t55);
and(z88, b88, r21);
and(a89, a88, r21);
and(b89, x88, u21, s21);
and(c89, y88, d15, s21);
and(d89, y88, f15, y21);
and(e89, x88, w21, y21);
and(f89, x88, q22, o22);
and(g89, y88, x15, o22);
and(h89, x88, u22, s22);
and(i89, y88, b16, s22);
and(j89, z4, k88, o88, s79, t81);
not(t_732, v87);
not(t_733, g70);
or(k89, t_732, t_733);
not(l89, x87);
and(m89, n88, o86);
not(n89, a88);
not(t_734, q70);
not(t_735, l88);
or(o89, t_734, t_735);
not(t_736, r70);
not(t_737, m88);
or(p89, t_736, t_737);
not(q89, b88);
not(r89, c88);
not(s89, d88);
not(t_738, i72);
not(t_739, c88);
or(t89, t_738, t_739);
not(t_740, j72);
not(t_741, d88);
or(u89, t_740, t_741);
not(t_742, h88);
not(t_743, a73);
or(v89, t_742, t_743);
not(t_744, g88);
not(t_745, b73);
or(w89, t_744, t_745);
not(t_746, s58);
not(t_747, x87);
or(x89, t_746, t_747);
not(y89, l88);
not(z89, m88);
and(a90, l77, n88);
or(b90, f30, v36, s87, r87);
or(c90, g30, w36, u87, t87);
or(d90, q87, b31, u77, p49);
or(e90, v37, i87, n49);
or(f90, x37, j87, m49);
or(g90, d38, k87, b60);
or(h90, e38, l87, u55);
and(i90, n89, p21, j21);
and(j90, q89, q21, l21);
and(k90, e90, u21, s21);
and(l90, f90, u21, s21);
and(m90, g90, d15, s21);
and(n90, h90, d15, s21);
and(o90, g90, f15, y21);
and(p90, h90, f15, y21);
and(q90, e90, w21, y21);
and(r90, f90, w21, y21);
and(s90, f90, q22, o22);
and(t90, e90, q22, o22);
and(u90, g90, x15, o22);
and(v90, h90, x15, o22);
and(w90, f90, u22, s22);
and(x90, e90, u22, s22);
and(y90, g90, b16, s22);
and(z90, h90, b16, s22);
not(t_748, w87);
not(t_749, k89);
or(a91, t_748, t_749);
not(t_750, y89);
not(t_751, w63);
or(b91, t_750, t_751);
not(t_752, z89);
not(t_753, y63);
or(c91, t_752, t_753);
not(t_754, r89);
not(t_755, d66);
or(d91, t_754, t_755);
not(t_756, s89);
not(t_757, e66);
or(e91, t_756, t_757);
not(t_758, i88);
not(t_759, v89);
or(f91, t_758, t_759);
not(t_760, j88);
not(t_761, w89);
or(g91, t_760, t_761);
not(t_762, l89);
not(t_763, q52);
or(h91, t_762, t_763);
or(i91, j30, a37, i89, h89);
or(j91, k30, z36, g89, f89);
not(k91, a91);
not(t_764, o89);
not(t_765, b91);
or(l91, t_764, t_765);
not(t_766, p89);
not(t_767, c91);
or(m91, t_766, t_767);
not(t_768, t89);
not(t_769, d91);
or(n91, t_768, t_769);
not(t_770, u89);
not(t_771, e91);
or(o91, t_770, t_771);
not(p91, f91);
not(q91, g91);
not(t_772, c73);
not(t_773, f91);
or(r91, t_772, t_773);
not(t_774, d73);
not(t_775, g91);
or(s91, t_774, t_775);
not(t_776, r58);
not(t_777, a91);
or(t91, t_776, t_777);
not(t_778, x89);
not(t_779, h91);
or(u91, t_778, t_779);
or(v91, l30, b37, v90, s90);
or(w91, m30, c37, z90, w90);
or(x91, n30, e37, y90, x90);
or(y91, o30, d37, u90, t90);
not(t_780, t69);
not(t_781, u91);
or(z91, t_780, t_781);
not(a92, l91);
not(b92, m91);
not(t_782, y70);
not(t_783, m91);
or(c92, t_782, t_783);
not(t_784, z70);
not(t_785, l91);
or(d92, t_784, t_785);
not(t_786, g71);
not(t_787, o91);
or(e92, t_786, t_787);
not(t_788, h71);
not(t_789, n91);
or(f92, t_788, t_789);
not(g92, n91);
not(h92, o91);
not(t_790, p91);
not(t_791, l67);
or(i92, t_790, t_791);
not(t_792, q91);
not(t_793, m67);
or(j92, t_792, t_793);
not(t_794, k91);
not(t_795, p52);
or(k92, t_794, t_795);
not(l92, u91);
not(t_796, l92);
not(t_797, w62);
or(m92, t_796, t_797);
not(t_798, b92);
not(t_799, m64);
or(n92, t_798, t_799);
not(t_800, a92);
not(t_801, n64);
or(o92, t_800, t_801);
not(t_802, h92);
not(t_803, y64);
or(p92, t_802, t_803);
not(t_804, g92);
not(t_805, b65);
or(q92, t_804, t_805);
not(t_806, r91);
not(t_807, i92);
or(r92, t_806, t_807);
not(t_808, s91);
not(t_809, j92);
or(s92, t_808, t_809);
not(t_810, t91);
not(t_811, k92);
or(t92, t_810, t_811);
not(t_812, z91);
not(t_813, m92);
or(u92, t_812, t_813);
not(t_814, u69);
not(t_815, t92);
or(v92, t_814, t_815);
not(t_816, c92);
not(t_817, n92);
or(w92, t_816, t_817);
not(t_818, d92);
not(t_819, o92);
or(x92, t_818, t_819);
not(t_820, e92);
not(t_821, p92);
or(y92, t_820, t_821);
not(t_822, f92);
not(t_823, q92);
or(z92, t_822, t_823);
not(t_824, n72);
not(t_825, s92);
or(a93, t_824, t_825);
not(t_826, o72);
not(t_827, r92);
or(b93, t_826, t_827);
not(c93, r92);
not(d93, s92);
not(e93, t92);
not(f93, u92);
not(t_828, e93);
not(t_829, x62);
or(g93, t_828, t_829);
not(t_830, k70);
not(t_831, u92);
or(h93, t_830, t_831);
not(i93, w92);
not(j93, x92);
not(k93, y92);
not(l93, z92);
not(t_832, w71);
not(t_833, z92);
or(m93, t_832, t_833);
not(t_834, x71);
not(t_835, y92);
or(n93, t_834, t_835);
not(t_836, d93);
not(t_837, o66);
or(o93, t_836, t_837);
not(t_838, c93);
not(t_839, r66);
or(p93, t_838, t_839);
not(t_840, j59);
not(t_841, x92);
or(q93, t_840, t_841);
not(t_842, k59);
not(t_843, w92);
or(r93, t_842, t_843);
not(t_844, v92);
not(t_845, g93);
or(s93, t_844, t_845);
not(t_846, f93);
not(t_847, t63);
or(t93, t_846, t_847);
not(t_848, l93);
not(t_849, p65);
or(u93, t_848, t_849);
not(t_850, k93);
not(t_851, q65);
or(v93, t_850, t_851);
not(t_852, a93);
not(t_853, o93);
or(w93, t_852, t_853);
not(t_854, b93);
not(t_855, p93);
or(x93, t_854, t_855);
not(t_856, j93);
not(t_857, b54);
or(y93, t_856, t_857);
not(t_858, i93);
not(t_859, c54);
or(z93, t_858, t_859);
not(a94, s93);
not(t_860, j70);
not(t_861, s93);
or(b94, t_860, t_861);
not(t_862, h93);
not(t_863, t93);
or(c94, t_862, t_863);
not(t_864, m93);
not(t_865, u93);
or(d94, t_864, t_865);
not(t_866, n93);
not(t_867, v93);
or(e94, t_866, t_867);
not(t_868, a72);
not(t_869, x93);
or(f94, t_868, t_869);
not(t_870, b72);
not(t_871, w93);
or(g94, t_870, t_871);
not(h94, w93);
not(i94, x93);
not(t_872, q93);
not(t_873, y93);
or(j94, t_872, t_873);
not(t_874, r93);
not(t_875, z93);
or(k94, t_874, t_875);
not(t_876, b70);
not(t_877, c94);
or(l94, t_876, t_877);
not(t_878, a94);
not(t_879, s63);
or(m94, t_878, t_879);
not(n94, c94);
not(t_880, k71);
not(t_881, e94);
or(o94, t_880, t_881);
not(t_882, l71);
not(t_883, d94);
or(p94, t_882, t_883);
not(q94, d94);
not(r94, e94);
not(t_884, i94);
not(t_885, s65);
or(s94, t_884, t_885);
not(t_886, h94);
not(t_887, t65);
or(t94, t_886, t_887);
not(t_888, e59);
not(t_889, k94);
or(u94, t_888, t_889);
not(t_890, f59);
not(t_891, j94);
or(v94, t_890, t_891);
not(w94, j94);
not(x94, k94);
not(t_892, n94);
not(t_893, k63);
or(y94, t_892, t_893);
not(t_894, b94);
not(t_895, m94);
or(z94, t_894, t_895);
not(t_896, r94);
not(t_897, g65);
or(a95, t_896, t_897);
not(t_898, q94);
not(t_899, h65);
or(b95, t_898, t_899);
not(t_900, f94);
not(t_901, s94);
or(c95, t_900, t_901);
not(t_902, g94);
not(t_903, t94);
or(d95, t_902, t_903);
not(t_904, x94);
not(t_905, r53);
or(e95, t_904, t_905);
not(t_906, w94);
not(t_907, s53);
or(f95, t_906, t_907);
not(t_908, a70);
not(t_909, z94);
or(g95, t_908, t_909);
not(t_910, l94);
not(t_911, y94);
or(h95, t_910, t_911);
not(i95, z94);
not(t_912, o94);
not(t_913, a95);
or(j95, t_912, t_913);
not(t_914, p94);
not(t_915, b95);
or(k95, t_914, t_915);
not(l95, c95);
not(m95, d95);
not(t_916, q72);
not(t_917, c95);
or(n95, t_916, t_917);
not(t_918, r72);
not(t_919, d95);
or(o95, t_918, t_919);
not(t_920, u94);
not(t_921, e95);
or(p95, t_920, t_921);
not(t_922, v94);
not(t_923, f95);
or(q95, t_922, t_923);
and(r95, q95, w74, t15);
and(s95, p95, l70, t15);
and(t95, p95, l81, f5);
and(u95, q95, o79, f5);
and(v95, k95, v75, c16);
and(w95, j95, d72, c16);
and(x95, j95, u80, a5);
and(y95, k95, t78, a5);
not(t_924, i95);
not(t_925, j63);
or(z95, t_924, t_925);
not(a96, h95);
not(t_926, o63);
not(t_927, h95);
or(b96, t_926, t_927);
not(t_928, l95);
not(t_929, y66);
or(c96, t_928, t_929);
not(t_930, m95);
not(t_931, z66);
or(d96, t_930, t_931);
or(e96, t95, u95, s95, r95);
or(f96, x95, y95, w95, v95);
not(t_932, g95);
not(t_933, z95);
or(g96, t_932, t_933);
not(t_934, a96);
not(t_935, o60);
or(h96, t_934, t_935);
not(t_936, n95);
not(t_937, c96);
or(i96, t_936, t_937);
not(t_938, o95);
not(t_939, d96);
or(j96, t_938, t_939);
not(k96, e96);
not(l96, f96);
not(m96, g96);
not(t_940, n63);
not(t_941, g96);
or(n96, t_940, t_941);
not(t_942, b96);
not(t_943, h96);
or(o96, t_942, t_943);
not(p96, i96);
not(q96, j96);
not(t_944, y72);
not(t_945, i96);
or(r96, t_944, t_945);
not(t_946, z72);
not(t_947, j96);
or(s96, t_946, t_947);
and(t96, f5, o96);
not(t_948, m96);
not(t_949, n60);
or(u96, t_948, t_949);
not(t_950, p96);
not(t_951, i67);
or(v96, t_950, t_951);
not(t_952, q96);
not(t_953, j67);
or(w96, t_952, t_953);
not(t_954, n96);
not(t_955, u96);
or(x96, t_954, t_955);
not(t_956, r96);
not(t_957, v96);
or(y96, t_956, t_957);
not(t_958, s96);
not(t_959, w96);
or(z96, t_958, t_959);
and(a97, a5, z96);
not(b97, x96);
not(c97, y96);
and(d97, b97, t15);
and(e97, c97, c16);
or(f97, t96, d97);
or(g97, a97, e97);
not(t_960, k96);
not(t_961, f97);
or(h97, t_960, t_961);
not(i97, f97);
not(t_962, l96);
not(t_963, g97);
or(j97, t_962, t_963);
not(k97, g97);
not(t_964, i97);
not(t_965, e96);
or(l97, t_964, t_965);
not(t_966, k97);
not(t_967, f96);
or(m97, t_966, t_967);
not(t_968, l97);
not(t_969, h97);
or(n97, t_968, t_969);
not(t_970, m97);
not(t_971, j97);
or(o97, t_970, t_971);
and(p97, n97, y14, j21);
and(q97, o97, z14, l21);
not(r97, n97);
not(s97, o97);
and(t97, r97, a15);
and(u97, s97, a15);
or(v97, u97, z88);
or(w97, t97, a89);
and(x97, v97, m21);
and(y97, v97, m21);
and(z97, w97, m21);
and(a98, w97, m21);
or(b98, g31, y97);
or(c98, h31, x97);
or(d98, i31, a98);
or(e98, j31, z97);
and(f98, d98, v21, t21);
and(g98, b98, e15, t21);
and(h98, b98, g15, z21);
and(i98, d98, x21, z21);
and(j98, e98, p22, n22);
and(k98, c98, w15, n22);
and(l98, e98, t22, r22);
and(m98, c98, a16, r22);
or(n98, d30, k37, m98, l98);
or(o98, e30, j37, k98, j98);
and(p98, n98, x30);
and(q98, o98, y30);
buf(w5, n1);
buf(x5, i3);
buf(y5, i5);
buf(z6, i32);
buf(a7, i32);
buf(b7, i32);
buf(c7, i32);
endmodule
module top;
	parameter in_width = 178,
		patterns = 5000,
		step = 1;
	reg [1:in_width] in_mem[1:patterns];
	integer index;

	wire i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,
		i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,
		i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,
		i30,i31,i32,i33,i34,i35,i36,i37,i38,i39,
		i40,i41,i42,i43,i44,i45,i46,i47,i48,i49,
		i50,i51,i52,i53,i54,i55,i56,i57,i58,i59,
		i60,i61,i62,i63,i64,i65,i66,i67,i68,i69,
		i70,i71,i72,i73,i74,i75,i76,i77,i78,i79,
		i80,i81,i82,i83,i84,i85,i86,i87,i88,i89,
		i90,i91,i92,i93,i94,i95,i96,i97,i98,i99,
		i100,i101,i102,i103,i104,i105,i106,i107,i108,i109,
		i110,i111,i112,i113,i114,i115,i116,i117,i118,i119,
		i120,i121,i122,i123,i124,i125,i126,i127,i128,i129,
		i130,i131,i132,i133,i134,i135,i136,i137,i138,i139,
		i140,i141,i142,i143,i144,i145,i146,i147,i148,i149,
		i150,i151,i152,i153,i154,i155,i156,i157,i158,i159,
		i160,i161,i162,i163,i164,i165,i166,i167,i168,i169,
		i170,i171,i172,i173,i174,i175,i176,i177;

	assign {i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,
		i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,
		i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,
		i30,i31,i32,i33,i34,i35,i36,i37,i38,i39,
		i40,i41,i42,i43,i44,i45,i46,i47,i48,i49,
		i50,i51,i52,i53,i54,i55,i56,i57,i58,i59,
		i60,i61,i62,i63,i64,i65,i66,i67,i68,i69,
		i70,i71,i72,i73,i74,i75,i76,i77,i78,i79,
		i80,i81,i82,i83,i84,i85,i86,i87,i88,i89,
		i90,i91,i92,i93,i94,i95,i96,i97,i98,i99,
		i100,i101,i102,i103,i104,i105,i106,i107,i108,i109,
		i110,i111,i112,i113,i114,i115,i116,i117,i118,i119,
		i120,i121,i122,i123,i124,i125,i126,i127,i128,i129,
		i130,i131,i132,i133,i134,i135,i136,i137,i138,i139,
		i140,i141,i142,i143,i144,i145,i146,i147,i148,i149,
		i150,i151,i152,i153,i154,i155,i156,i157,i158,i159,
		i160,i161,i162,i163,i164,i165,i166,i167,i168,i169,
		i170,i171,i172,i173,i174,i175,i176,i177} = 
		$getpattern(in_mem[index]);

	initial $monitor($time,,o0,o1,o2,o3,o4,o5,o6,o7,o8,o9,
		o10,o11,o12,o13,o14,o15,o16,o17,o18,o19,
		o20,o21,o22,o23,o24,o25,o26,o27,o28,o29,
		o30,o31,o32,o33,o34,o35,o36,o37,o38,o39,
		o40,o41,o42,o43,o44,o45,o46,o47,o48,o49,
		o50,o51,o52,o53,o54,o55,o56,o57,o58,o59,
		o60,o61,o62,o63,o64,o65,o66,o67,o68,o69,
		o70,o71,o72,o73,o74,o75,o76,o77,o78,o79,
		o80,o81,o82,o83,o84,o85,o86,o87,o88,o89,
		o90,o91,o92,o93,o94,o95,o96,o97,o98,o99,
		o100,o101,o102,o103,o104,o105,o106,o107,o108,o109,
		o110,o111,o112,o113,o114,o115,o116,o117,o118,o119,
		o120,o121,o122);
	initial
		begin
			$readmemb("patt.mem", in_mem);
			for(index = 1; index <= patterns; index = index + 1)
				#step;
		end

	foobar cct(o0,o1,o2,o3,o4,o5,o6,o7,o8,o9,
		o10,o11,o12,o13,o14,o15,o16,o17,o18,o19,
		o20,o21,o22,o23,o24,o25,o26,o27,o28,o29,
		o30,o31,o32,o33,o34,o35,o36,o37,o38,o39,
		o40,o41,o42,o43,o44,o45,o46,o47,o48,o49,
		o50,o51,o52,o53,o54,o55,o56,o57,o58,o59,
		o60,o61,o62,o63,o64,o65,o66,o67,o68,o69,
		o70,o71,o72,o73,o74,o75,o76,o77,o78,o79,
		o80,o81,o82,o83,o84,o85,o86,o87,o88,o89,
		o90,o91,o92,o93,o94,o95,o96,o97,o98,o99,
		o100,o101,o102,o103,o104,o105,o106,o107,o108,o109,
		o110,o111,o112,o113,o114,o115,o116,o117,o118,o119,
		o120,o121,o122,i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,
		i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,
		i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,
		i30,i31,i32,i33,i34,i35,i36,i37,i38,i39,
		i40,i41,i42,i43,i44,i45,i46,i47,i48,i49,
		i50,i51,i52,i53,i54,i55,i56,i57,i58,i59,
		i60,i61,i62,i63,i64,i65,i66,i67,i68,i69,
		i70,i71,i72,i73,i74,i75,i76,i77,i78,i79,
		i80,i81,i82,i83,i84,i85,i86,i87,i88,i89,
		i90,i91,i92,i93,i94,i95,i96,i97,i98,i99,
		i100,i101,i102,i103,i104,i105,i106,i107,i108,i109,
		i110,i111,i112,i113,i114,i115,i116,i117,i118,i119,
		i120,i121,i122,i123,i124,i125,i126,i127,i128,i129,
		i130,i131,i132,i133,i134,i135,i136,i137,i138,i139,
		i140,i141,i142,i143,i144,i145,i146,i147,i148,i149,
		i150,i151,i152,i153,i154,i155,i156,i157,i158,i159,
		i160,i161,i162,i163,i164,i165,i166,i167,i168,i169,
		i170,i171,i172,i173,i174,i175,i176,i177);
endmodule
