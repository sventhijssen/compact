module s444(VDD,CK,G0,G1,G107,G108,G118,G119,G167,G168,G2);
input VDD,CK,G0,G1,G2;
output G118,G167,G107,G119,G168,G108;

  wire G11,G37,G12,G41,G13,G45,G14,G49,G15,G58,G16,G62,G17,G66,G18,G70,G19,G80,
    G20,G84,G21,G88,G22,G92,G23,G101,G24,G162BF,G25,G109,G26,G110,G27,G111,G28,
    G112,G29,G113,G30,G114,G31,G155,IIII372,IIII382,IIII318,G34,IIII180,G35,
    G77,G135,G36,G78,G144,G32,G74,G142,IIII392,G55,G102,G136,G156,G56,G143,
    G161,IIII321,G53,IIII324,G76,G150,IIII336,G152,G160,G106,G43,IIII182,G99,
    G139,G153,G157,G103,G38,G40,G60,G57,G79,G97,G42,G44,G46,G48,IIII105,G162,
    G166,G50,G52,G82,G59,G61,G63,G65,G67,G69,G71,G73,G81,G83,G85,G87,G89,G91,
    G94,G96,G122,G121,G124,G125,G126,G127,G154,G158,G159,G100,G104,G105,G115,
    G117,G163,G165,G116,G164,G141,G137,G138,G140,G133,G134,G145,G146,G147,G131,
    G129,IIII181,IIII190,IIII200,G47,IIII210,G51,G120,G128,G132,G123,G151,
    IIII191,IIII192,IIII201,IIII202,G149,G130,IIII211,IIII212,G148,IIII225,
    IIII235,G64,IIII245,G68,IIII255,G72,IIII226,IIII227,IIII236,IIII237,
    IIII246,IIII247,IIII256,IIII257,IIII271,IIII281,G86,IIII291,G90,IIII302,
    G95,IIII272,IIII273,IIII282,IIII283,IIII292,IIII293,IIII303,IIII304,G33,
    G54,G75,G98,G93;

  FD1 DFF_0(CK,G11,G37);
  FD1 DFF_1(CK,G12,G41);
  FD1 DFF_2(CK,G13,G45);
  FD1 DFF_3(CK,G14,G49);
  FD1 DFF_4(CK,G15,G58);
  FD1 DFF_5(CK,G16,G62);
  FD1 DFF_6(CK,G17,G66);
  FD1 DFF_7(CK,G18,G70);
  FD1 DFF_8(CK,G19,G80);
  FD1 DFF_9(CK,G20,G84);
  FD1 DFF_10(CK,G21,G88);
  FD1 DFF_11(CK,G22,G92);
  FD1 DFF_12(CK,G23,G101);
  FD1 DFF_13(CK,G24,G162BF);
  FD1 DFF_14(CK,G25,G109);
  FD1 DFF_15(CK,G26,G110);
  FD1 DFF_16(CK,G27,G111);
  FD1 DFF_17(CK,G28,G112);
  FD1 DFF_18(CK,G29,G113);
  FD1 DFF_19(CK,G30,G114);
  FD1 DFF_20(CK,G31,G155);
  IV  NOT_0(IIII372,G0);
  IV  NOT_1(IIII382,G1);
  IV  NOT_2(IIII318,G2);
  IV  NOT_3(G34,G11);
  IV  NOT_4(IIII180,G11);
  IV  NOT_5(G35,G12);
  IV  NOT_6(G77,G20);
  IV  NOT_7(G135,G20);
  IV  NOT_8(G36,G13);
  IV  NOT_9(G78,G21);
  IV  NOT_10(G144,G21);
  IV  NOT_11(G32,G14);
  IV  NOT_12(G74,G22);
  IV  NOT_13(G142,G22);
  IV  NOT_14(IIII392,G30);
  IV  NOT_15(G55,G15);
  IV  NOT_16(G102,G23);
  IV  NOT_17(G136,G23);
  IV  NOT_18(G156,G31);
  IV  NOT_19(G56,G16);
  IV  NOT_20(G143,G24);
  IV  NOT_21(G161,G17);
  IV  NOT_22(IIII321,G25);
  IV  NOT_23(G53,G18);
  IV  NOT_24(IIII324,G26);
  IV  NOT_25(G76,G19);
  IV  NOT_26(G150,G19);
  IV  NOT_27(IIII336,G27);
  IV  NOT_28(G119,G28);
  IV  NOT_29(G167,G29);
  IV  NOT_30(G152,IIII372);
  IV  NOT_31(G160,IIII382);
  IV  NOT_32(G106,IIII318);
  IV  NOT_33(G43,G34);
  IV  NOT_34(IIII182,IIII180);
  IV  NOT_35(G168,IIII392);
  IV  NOT_36(G107,IIII321);
  IV  NOT_37(G108,IIII324);
  IV  NOT_38(G118,IIII336);
  IV  NOT_39(G99,G152);
  IV  NOT_40(G139,G152);
  IV  NOT_41(G153,G152);
  IV  NOT_42(G157,G160);
  IV  NOT_43(G103,G106);
  IV  NOT_44(G38,G40);
  IV  NOT_45(G60,G57);
  IV  NOT_46(G79,G97);
  IV  NOT_47(G42,G44);
  IV  NOT_48(G46,G48);
  IV  NOT_49(IIII105,G162);
  IV  NOT_50(G166,G162);
  IV  NOT_51(G50,G52);
  IV  NOT_52(G82,G79);
  IV  NOT_53(G162BF,IIII105);
  IV  NOT_54(G59,G61);
  IV  NOT_55(G63,G65);
  IV  NOT_56(G67,G69);
  IV  NOT_57(G71,G73);
  IV  NOT_58(G81,G83);
  IV  NOT_59(G85,G87);
  IV  NOT_60(G89,G91);
  IV  NOT_61(G94,G96);
  AN2 AND2_0(G122,G24,G121);
  AN3 AND3_0(G124,G139,G22,G150);
  AN3 AND3_1(G125,G139,G20,G19);
  AN2 AND2_1(G126,G139,G21);
  AN2 AND2_2(G127,G139,G24);
  AN2 AND2_3(G154,G158,G159);
  AN2 AND2_4(G100,G104,G105);
  AN2 AND2_5(G155,G154,G153);
  AN2 AND2_6(G101,G100,G99);
  AN3 AND3_2(G115,G161,G117,G162);
  AN3 AND3_3(G163,G161,G165,G162);
  AN2 AND2_7(G116,G117,G166);
  AN2 AND2_8(G164,G165,G166);
  OR3 OR3_0(G141,G24,G22,G21);
  OR3 OR3_1(G137,G136,G20,G19);
  OR2 OR2_0(G138,G136,G142);
  OR4 OR4_0(G140,G24,G21,G20,G150);
  OR4 OR4_1(G133,G152,G136,G22,G144);
  OR3 OR3_2(G134,G152,G142,G21);
  OR4 OR4_2(G145,G152,G142,G20,G19);
  OR2 OR2_1(G146,G152,G143);
  OR2 OR2_2(G147,G152,G144);
  OR2 OR2_3(G158,G31,G160);
  OR2 OR2_4(G104,G23,G106);
  OR4 OR4_3(G131,G144,G22,G23,G129);
  OR2 OR2_5(G159,G156,G157);
  OR2 OR2_6(G105,G102,G103);
  ND2 NAND2_0(IIII181,G11,IIII180);
  ND2 NAND2_1(G129,G19,G135);
  ND4 NAND4_0(G121,G19,G135,G142,G136);
  ND2 NAND2_2(IIII190,G12,G43);
  ND2 NAND2_3(G40,IIII181,IIII182);
  ND2 NAND2_4(IIII200,G13,G47);
  ND2 NAND2_5(IIII210,G14,G51);
  ND2 NAND2_6(G120,G150,G128);
  ND2 NAND2_7(G132,G133,G134);
  ND3 NAND3_0(G111,G140,G141,G139);
  ND4 NAND4_1(G123,G137,G138,G21,G139);
  ND4 NAND4_2(G151,G20,G144,G143,G139);
  ND3 NAND3_1(G117,G145,G146,G147);
  ND2 NAND2_8(IIII191,G12,IIII190);
  ND2 NAND2_9(IIII192,G43,IIII190);
  ND2 NAND2_10(IIII201,G13,IIII200);
  ND2 NAND2_11(IIII202,G47,IIII200);
  ND2 NAND2_12(G149,G131,G130);
  ND2 NAND2_13(IIII211,G14,IIII210);
  ND2 NAND2_14(IIII212,G51,IIII210);
  ND3 NAND3_2(G148,G150,G135,G132);
  ND2 NAND2_15(G44,IIII191,IIII192);
  ND2 NAND2_16(G48,IIII201,IIII202);
  ND2 NAND2_17(G162,G120,G149);
  ND2 NAND2_18(G52,IIII211,IIII212);
  ND2 NAND2_19(IIII225,G15,G60);
  ND2 NAND2_20(IIII235,G16,G64);
  ND2 NAND2_21(IIII245,G17,G68);
  ND2 NAND2_22(IIII255,G18,G72);
  ND2 NAND2_23(G165,G148,G149);
  ND2 NAND2_24(IIII226,G15,IIII225);
  ND2 NAND2_25(IIII227,G60,IIII225);
  ND2 NAND2_26(IIII236,G16,IIII235);
  ND2 NAND2_27(IIII237,G64,IIII235);
  ND2 NAND2_28(IIII246,G17,IIII245);
  ND2 NAND2_29(IIII247,G68,IIII245);
  ND2 NAND2_30(IIII256,G18,IIII255);
  ND2 NAND2_31(IIII257,G72,IIII255);
  ND2 NAND2_32(G61,IIII226,IIII227);
  ND2 NAND2_33(G65,IIII236,IIII237);
  ND2 NAND2_34(G69,IIII246,IIII247);
  ND2 NAND2_35(G73,IIII256,IIII257);
  ND2 NAND2_36(IIII271,G19,G82);
  ND2 NAND2_37(IIII281,G20,G86);
  ND2 NAND2_38(IIII291,G21,G90);
  ND2 NAND2_39(IIII302,G22,G95);
  ND2 NAND2_40(IIII272,G19,IIII271);
  ND2 NAND2_41(IIII273,G82,IIII271);
  ND2 NAND2_42(IIII282,G20,IIII281);
  ND2 NAND2_43(IIII283,G86,IIII281);
  ND2 NAND2_44(IIII292,G21,IIII291);
  ND2 NAND2_45(IIII293,G90,IIII291);
  ND2 NAND2_46(IIII303,G22,IIII302);
  ND2 NAND2_47(IIII304,G95,IIII302);
  ND2 NAND2_48(G83,IIII272,IIII273);
  ND2 NAND2_49(G87,IIII282,IIII283);
  ND2 NAND2_50(G91,IIII292,IIII293);
  ND2 NAND2_51(G96,IIII303,IIII304);
  NR3 NOR3_0(G33,G11,G12,G13);
  NR3 NOR3_1(G54,G15,G16,G17);
  NR3 NOR3_2(G75,G19,G20,G21);
  NR2 NOR2_0(G47,G34,G35);
  NR3 NOR3_3(G51,G34,G35,G36);
  NR2 NOR2_1(G98,G32,G33);
  NR4 NOR4_0(G128,G20,G144,G136,G152);
  NR2 NOR2_2(G130,G143,G152);
  NR2 NOR2_3(G57,G31,G98);
  NR2 NOR2_4(G64,G55,G57);
  NR3 NOR3_4(G68,G55,G56,G57);
  NR4 NOR4_1(G72,G55,G56,G161,G57);
  NR3 NOR3_5(G97,G53,G57,G54);
  NR2 NOR2_5(G109,G122,G123);
  NR4 NOR4_2(G110,G124,G125,G126,G127);
  NR2 NOR2_6(G114,G150,G151);
  NR3 NOR3_6(G37,G98,G38,G152);
  NR2 NOR2_7(G86,G76,G79);
  NR3 NOR3_7(G90,G76,G77,G79);
  NR3 NOR3_8(G93,G74,G79,G75);
  NR4 NOR4_3(G95,G76,G77,G78,G79);
  NR3 NOR3_9(G41,G98,G42,G152);
  NR3 NOR3_10(G45,G98,G46,G152);
  NR3 NOR3_11(G49,G98,G50,G152);
  NR2 NOR2_8(G112,G115,G116);
  NR2 NOR2_9(G113,G163,G164);
  NR3 NOR3_12(G58,G97,G59,G152);
  NR3 NOR3_13(G62,G97,G63,G152);
  NR3 NOR3_14(G66,G97,G67,G152);
  NR3 NOR3_15(G70,G97,G71,G152);
  NR3 NOR3_16(G80,G93,G81,G152);
  NR3 NOR3_17(G84,G93,G85,G152);
  NR3 NOR3_18(G88,G93,G89,G152);
  NR3 NOR3_19(G92,G93,G94,G152);

endmodule
