// IWLS benchmark module "pair" printed on Wed May 29 16:09:22 2002
module pair(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2, b2, c2, d2, e2, f2, g2, h2, i2, j2, k2, l2, m2, n2, o2, p2, q2, r2, s2, t2, u2, v2, w2, x2, y2, z2, a3, b3, c3, d3, e3, f3, g3, h3, i3, j3, k3, l3, m3, n3, o3, p3, q3, r3, s3, t3, u3, v3, w3, x3, y3, z3, a4, b4, c4, d4, e4, f4, g4, h4, i4, j4, k4, l4, m4, n4, o4, p4, q4, r4, s4, t4, u4, v4, w4, x4, y4, z4, a5, b5, c5, d5, e5, f5, g5, h5, i5, j5, k5, l5, m5, n5, o5, p5, q5, r5, s5, t5, u5, v5, w5, x5, y5, z5, a6, b6, c6, d6, e6, f6, g6, h6, i6, j6, k6, l6, m6, n6, o6, p6, q6, r6, s6, t6, u6, v6, w6, x6, y6, z6, a7, b7, c7, d7, e7, f7, g7, h7, i7, j7, k7, l7, m7, n7, o7, p7, q7, r7, s7, t7, u7, v7, w7, x7, y7, z7, a8, b8, c8, d8, e8, f8, g8, h8, i8, j8, k8, l8, m8, n8, o8, p8, q8, r8, s8, t8, u8, v8, w8, x8, y8, z8, a9, b9, c9, d9, e9, f9, g9, h9, i9, j9, k9, l9, m9, n9, o9, p9, q9, r9, s9, t9, u9, v9, w9, x9, y9, z9, a10, b10, c10, d10, e10, f10, g10, h10, i10, j10, k10, l10, m10, n10, o10, p10, q10, r10, s10, t10, u10, v10, w10, x10, y10);
input
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  t,
  u,
  v,
  w,
  y,
  z,
  a0,
  a1,
  a2,
  a3,
  a4,
  a5,
  b0,
  b1,
  b2,
  b3,
  b4,
  b5,
  c0,
  c1,
  c2,
  c3,
  c4,
  c5,
  d0,
  d1,
  d2,
  d3,
  d4,
  d5,
  e0,
  e1,
  e2,
  e3,
  e4,
  e5,
  f0,
  f1,
  f2,
  f3,
  f4,
  f5,
  g0,
  g1,
  g2,
  g3,
  g4,
  g5,
  h0,
  h1,
  h2,
  h3,
  h4,
  h5,
  i0,
  i1,
  i2,
  i3,
  i4,
  i5,
  j0,
  j1,
  j2,
  j3,
  j4,
  j5,
  k0,
  k1,
  k2,
  k3,
  k4,
  k5,
  l0,
  l1,
  l2,
  l3,
  l4,
  l5,
  m0,
  m1,
  m2,
  m3,
  m4,
  m5,
  n0,
  n1,
  n2,
  n3,
  n4,
  n5,
  o0,
  o1,
  o2,
  o3,
  o4,
  o5,
  p0,
  p1,
  p2,
  p3,
  p4,
  p5,
  q0,
  q1,
  q2,
  q3,
  q4,
  q5,
  r0,
  r1,
  r2,
  r3,
  r4,
  r5,
  s0,
  s1,
  s2,
  s3,
  s4,
  t0,
  t1,
  t2,
  t3,
  t4,
  u0,
  u1,
  u2,
  u3,
  u4,
  v0,
  v1,
  v2,
  v3,
  v4,
  w0,
  w1,
  w2,
  w3,
  w4,
  x0,
  x1,
  x2,
  x3,
  x4,
  y0,
  y1,
  y2,
  y3,
  y4,
  z0,
  z1,
  z2,
  z3,
  z4;
output
  h10,
  x10,
  i10,
  y10,
  j10,
  k10,
  l10,
  m10,
  n10,
  a6,
  a7,
  a8,
  a9,
  b6,
  b7,
  b8,
  b9,
  c6,
  c7,
  c8,
  c9,
  d6,
  d7,
  d8,
  d9,
  e6,
  e7,
  e8,
  e9,
  f6,
  f7,
  f8,
  f9,
  g6,
  g7,
  g8,
  g9,
  h6,
  h7,
  h8,
  h9,
  i6,
  i7,
  i8,
  i9,
  j6,
  j7,
  j8,
  j9,
  k6,
  k7,
  k8,
  k9,
  l6,
  l7,
  l8,
  l9,
  m6,
  m7,
  m8,
  m9,
  n6,
  n7,
  n8,
  n9,
  o10,
  o6,
  o7,
  o8,
  o9,
  p6,
  p7,
  p8,
  p9,
  q6,
  q7,
  q8,
  q9,
  r6,
  r7,
  r8,
  r9,
  s5,
  s6,
  s7,
  s8,
  s9,
  t5,
  t6,
  t7,
  t8,
  t9,
  u5,
  u6,
  u7,
  u8,
  u9,
  v5,
  v6,
  v7,
  v8,
  v9,
  w5,
  w6,
  w7,
  w8,
  w9,
  x5,
  x6,
  x7,
  x8,
  x9,
  y5,
  y6,
  y7,
  y8,
  y9,
  z5,
  z6,
  z7,
  z8,
  z9,
  p10,
  a10,
  q10,
  b10,
  r10,
  c10,
  s10,
  d10,
  t10,
  e10,
  u10,
  f10,
  v10,
  g10,
  w10;
wire
  w39,
  \[77] ,
  \[78] ,
  w53,
  \[79] ,
  h20,
  h22,
  h31,
  h32,
  h40,
  \[80] ,
  \[81] ,
  \[82] ,
  \[83] ,
  \[84] ,
  \[85] ,
  x23,
  x29,
  \[86] ,
  \[87] ,
  \[88] ,
  x53,
  \[89] ,
  i19,
  i33,
  i44,
  \[90] ,
  \[91] ,
  \[92] ,
  \[93] ,
  \[94] ,
  y18,
  \[95] ,
  \[96] ,
  \[97] ,
  \[100] ,
  y43,
  y47,
  y48,
  \[98] ,
  y50,
  \[101] ,
  \[99] ,
  \[102] ,
  j18,
  \[103] ,
  j26,
  j27,
  \[104] ,
  \[105] ,
  j47,
  j50,
  j51,
  \[106] ,
  \[107] ,
  \[108] ,
  \[0] ,
  \[109] ,
  \[1] ,
  \[2] ,
  \[200] ,
  \[3] ,
  \[201] ,
  \[4] ,
  \[202] ,
  \[5] ,
  z22,
  \[203] ,
  \[6] ,
  z30,
  \[204] ,
  \[7] ,
  z40,
  \[110] ,
  \[205] ,
  \[8] ,
  z50,
  \[111] ,
  \[206] ,
  \[9] ,
  \[112] ,
  k20,
  \[113] ,
  \[114] ,
  \[209] ,
  k40,
  \[115] ,
  k45,
  \[116] ,
  \[117] ,
  \[118] ,
  \[210] ,
  \[211] ,
  \[212] ,
  \[121] ,
  \[122] ,
  \[123] ,
  \[124] ,
  l37,
  \[125] ,
  l51,
  \[126] ,
  \[128] ,
  \[129] ,
  \[130] ,
  \[131] ,
  \[132] ,
  m16,
  m19,
  \[133] ,
  \[134] ,
  \[135] ,
  m53,
  \[136] ,
  \[231] ,
  \[232] ,
  \[143] ,
  \[144] ,
  \[239] ,
  n38,
  n40,
  n43,
  \[145] ,
  n44,
  n50,
  \[146] ,
  \[241] ,
  \[243] ,
  \[247] ,
  o26,
  \[249] ,
  \[155] ,
  o49,
  \[156] ,
  \[157] ,
  \[158] ,
  \[159] ,
  \[252] ,
  \[253] ,
  \[254] ,
  \[160] ,
  \[255] ,
  \[256] ,
  \[257] ,
  p21,
  p22,
  \[163] ,
  p25,
  \[258] ,
  \[164] ,
  p36,
  \[259] ,
  \[165] ,
  p47,
  \[166] ,
  \[167] ,
  a26,
  \[168] ,
  a28,
  \[169] ,
  \[260] ,
  \[261] ,
  \[262] ,
  \[10] ,
  \[263] ,
  \[11] ,
  \[12] ,
  \[170] ,
  \[13] ,
  \[171] ,
  \[14] ,
  \[172] ,
  q19,
  \[15] ,
  \[173] ,
  \[16] ,
  \[174] ,
  q39,
  \[17] ,
  q42,
  \[175] ,
  \[18] ,
  \[176] ,
  \[177] ,
  b17,
  b18,
  \[178] ,
  b32,
  \[179] ,
  b46,
  \[21] ,
  \[22] ,
  \[180] ,
  \[23] ,
  \[181] ,
  \[24] ,
  \[182] ,
  r18,
  r20,
  \[183] ,
  \[26] ,
  \[184] ,
  r36,
  r38,
  \[27] ,
  \[185] ,
  \[28] ,
  r50,
  \[186] ,
  \[29] ,
  \[187] ,
  c25,
  \[188] ,
  \[189] ,
  c52,
  c54,
  \[30] ,
  \[31] ,
  \[32] ,
  \[190] ,
  \[33] ,
  \[191] ,
  \[34] ,
  s16,
  \[35] ,
  \[193] ,
  s24,
  \[36] ,
  \[194] ,
  \[37] ,
  \[195] ,
  \[38] ,
  \[39] ,
  \[197] ,
  d21,
  \[198] ,
  d31,
  \[199] ,
  \[40] ,
  \[41] ,
  \[42] ,
  \[43] ,
  \[44] ,
  \[45] ,
  t20,
  t22,
  \[46] ,
  \[47] ,
  \[48] ,
  \[49] ,
  e19,
  e29,
  e52,
  \[50] ,
  \[51] ,
  \[52] ,
  \[53] ,
  \[54] ,
  u19,
  \[55] ,
  u22,
  \[56] ,
  \[57] ,
  \[58] ,
  u53,
  \[59] ,
  f50,
  \[60] ,
  \[61] ,
  \[62] ,
  \[63] ,
  \[64] ,
  v19,
  \[65] ,
  \[66] ,
  v38,
  \[67] ,
  v41,
  v42,
  v49,
  \[68] ,
  v50,
  \[69] ,
  g29,
  g41,
  g49,
  \[70] ,
  \[71] ,
  \[72] ,
  \[73] ,
  \[74] ,
  \[75] ,
  \[76] ,
  w32;
assign
  w39 = (q39 & (~j50 & p3)) | ((q39 & (j50 & ~p3)) | (n38 & h0)),
  \[77]  = e52 & (o3 & (n3 & (m3 & l3))),
  \[78]  = (~n38 & (e52 & l3)) | (n38 & (e52 & ~l3)),
  w53 = (\[187]  & ~c0) | (~l5 & ~c0),
  h10 = y,
  \[79]  = (~r38 & (e52 & m3)) | (r38 & (e52 & ~m3)),
  h20 = \[257]  & ~b18,
  h22 = \[231]  | ~t20,
  h31 = (\[261]  & (x2 & w2)) | (\[260]  & (~x2 & ~w2)),
  h32 = (b32 & (~e19 & a3)) | ((b32 & (e19 & ~a3)) | (z30 & j)),
  h40 = ~t3 & (~s3 & (~r3 & (~q3 & (~p3 & (~o3 & n3))))),
  \[80]  = (~v38 & (e52 & n3)) | (v38 & (e52 & ~n3)),
  \[81]  = (r38 & (~j50 & (~o3 & (n3 & m3)))) | ((r38 & (j50 & (\[79]  & (~o3 & ~n3)))) | ((j50 & (e52 & (~\[79]  & o3))) | ((~r38 & (e52 & o3)) | ((~j50 & (o3 & ~n3)) | ((\[79]  & (o3 & n3)) | \[175] ))))),
  \[82]  = (~q39 & (e52 & p3)) | ((q39 & (e52 & ~p3)) | \[175] ),
  \[83]  = (~w39 & (e52 & q3)) | ((w39 & (e52 & ~q3)) | \[175] ),
  \[84]  = (~n40 & (e52 & r3)) | (n40 & (e52 & ~r3)),
  x10 = \[135] ,
  \[85]  = (~z40 & (n40 & (~j50 & r3))) | ((~z40 & (e52 & (~\[84]  & s3))) | ((~z40 & (~j50 & s3)) | ((~n40 & (e52 & s3)) | ((z40 & \[84] ) | \[175] )))),
  x23 = (~d21 & (~v19 & s1)) | (~d21 & (v19 & ~s1)),
  x29 = (~\[172]  & (r20 & ~e19)) | ((~\[171]  & (r20 & e19)) | (~\[143]  & (r20 & q1))),
  \[86]  = (~z40 & (e52 & t3)) | ((z40 & (e52 & ~t3)) | \[175] ),
  \[87]  = (\[155]  & (~g41 & ~u3)) | ((\[155]  & (g41 & u3)) | (\[210]  & l3)),
  \[88]  = (\[155]  & (~v41 & v3)) | ((\[155]  & (v41 & ~v3)) | (\[210]  & m3)),
  x53 = (\[187]  & ~b0) | (m5 & ~b0),
  i10 = a5,
  \[89]  = (~\[198]  & (\[155]  & ~w3)) | ((\[198]  & (\[155]  & w3)) | (\[210]  & n3)),
  i19 = ~c1 & (~b1 & (~a1 & m19)),
  i33 = (w32 & (e19 & (~d3 & ~c3))) | (~\[190]  & (w32 & ~e19)),
  i44 = (~\[194]  & f4) | (q5 & ~j0),
  \[90]  = (~q42 & (l51 & x3)) | ((\[254]  & l51) | ((~l51 & o3) | z)),
  \[91]  = (~v42 & (l51 & y3)) | ((v42 & (l51 & ~y3)) | ((~l51 & p3) | z)),
  \[92]  = (~\[204]  & (l51 & ~z3)) | ((\[204]  & (l51 & z3)) | ((~l51 & q3) | z)),
  \[93]  = (\[155]  & (~n43 & a4)) | ((\[155]  & (n43 & ~a4)) | (\[210]  & r3)),
  \[94]  = (~y43 & (n43 & (~z50 & (l51 & a4)))) | ((\[182]  & (~y43 & (l51 & b4))) | ((y43 & (z50 & l51)) | ((~n43 & (l51 & b4)) | ((~l51 & s3) | z)))),
  y10 = \[136] ,
  y18 = \[164]  | r18,
  \[95]  = (~y43 & (l51 & c4)) | ((y43 & (l51 & ~c4)) | ((~l51 & t3) | z)),
  \[96]  = z | ~d4,
  \[97]  = (~e4 & d4) | ((e4 & ~d4) | z),
  \[100]  = (~v50 & (~n44 & ~h4)) | ((\[212]  & h4) | ((v50 & v3) | z)),
  y43 = (n43 & (~z50 & (b4 & a4))) | (~\[182]  & (n43 & ~b4)),
  y47 = \[185]  | (~y4 | (~x4 | ~w4)),
  y48 = (n5 & (~m5 & l5)) | z,
  \[98]  = (~\[194]  & ~f4) | ((\[194]  & f4) | z),
  y50 = (~m53 & r5) | \[160] ,
  \[101]  = (~i44 & i4) | ((i44 & ~i4) | z),
  j10 = \[121] ,
  \[99]  = (~\[243]  & \[212] ) | ((\[212]  & \[183] ) | ((\[212]  & g4) | ((v50 & u3) | z))),
  \[102]  = (~\[168]  & (~v50 & ~j4)) | ((\[168]  & (~v50 & j4)) | ((v50 & w3) | z)),
  j18 = (~\[164]  & (y18 & ~i1)) | h1,
  \[103]  = (~\[168]  & (~k45 & (~v50 & j4))) | ((~k45 & (~v50 & k4)) | ((v50 & x3) | z)),
  j26 = (~\[193]  & d2) | (q1 & ~l),
  j27 = ~\[166]  & (i2 & h2),
  \[104]  = (~k45 & (~v50 & l4)) | ((k45 & (~v50 & ~l4)) | ((v50 & y3) | z)),
  \[105]  = (\[169]  & (~b46 & ~v50)) | ((~b46 & (~v50 & m4)) | ((v50 & z3) | z)),
  j47 = ~\[184]  & (u4 & (t4 & s4)),
  j50 = (~\[146]  & ~e0) | (u53 & ~e0),
  j51 = ~y48 & (~m5 & l5),
  \[106]  = (~b46 & (~v50 & n4)) | ((b46 & (~v50 & ~n4)) | ((v50 & a4) | z)),
  \[107]  = (~\[158]  & (~v50 & ~o4)) | ((\[158]  & (~v50 & o4)) | ((v50 & b4) | z)),
  \[108]  = (~v50 & (q4 & (o4 & (n4 & (m4 & (l4 & (k4 & (j4 & h4)))))))) | (q4 & (o4 & (n4 & (m4 & (l4 & (k4 & (j4 & (h4 & z)))))))),
  \[0]  = (e3 & m) | ((a3 & n) | ((t2 & o) | ((o2 & s) | ((j2 & t) | ((g2 & u) | ((a2 & p) | ((x1 & q) | ((u1 & r) | ((d1 & v) | (y0 & w)))))))))),
  \[109]  = (~\[206]  & (~v50 & ~q4)) | ((\[206]  & (~v50 & q4)) | ((v50 & c4) | z)),
  \[1]  = (d3 & m) | ((z2 & n) | ((s2 & o) | ((m2 & s) | ((i2 & t) | ((d2 & u) | ((z1 & p) | ((w1 & q) | ((t1 & r) | ((c1 & v) | (x0 & w)))))))))),
  \[2]  = (c3 & m) | ((y2 & n) | ((r2 & o) | ((l2 & s) | ((h2 & t) | ((c2 & u) | ((y1 & p) | ((v1 & q) | ((s1 & r) | ((b1 & v) | (w0 & w)))))))))),
  \[200]  = (~e19 & ~q2) | ((e19 & q2) | ~r20),
  \[3]  = (b3 & m) | ((x2 & n) | ((q2 & o) | ((k2 & s) | ((f2 & t) | ((b2 & u) | ((r1 & q) | ((p1 & p) | ((m1 & r) | ((a1 & v) | (v0 & w)))))))))),
  \[201]  = (g29 & ~e19) | ((e29 & e19) | ~r20),
  \[4]  = (~\[249]  & o) | ((~\[181]  & s) | ((p21 & m) | ((~r20 & u) | ((~t20 & q) | ((w2 & n) | ((e2 & t) | ((q1 & p) | ((n1 & r) | ((l1 & w) | (z0 & v)))))))))),
  \[202]  = (~j50 & ~f3) | ((j50 & f3) | ~c52),
  \[5]  = (z4 & t0) | ((u4 & u0) | ((q4 & q0) | ((l4 & r0) | ((i4 & s0) | ((c4 & n0) | ((z3 & o0) | ((w3 & p0) | ((t3 & k0) | ((p3 & l0) | (i3 & m0)))))))))),
  z22 = (~r1 & (~q1 & ~b)) | ((~r1 & (~p1 & ~b)) | (~q1 & (~p1 & ~b))),
  \[203]  = (r36 & ~j50) | ((p36 & j50) | ~c52),
  \[6]  = (y4 & t0) | ((t4 & u0) | ((o4 & q0) | ((k4 & r0) | ((f4 & s0) | ((b4 & n0) | ((y3 & o0) | ((v3 & p0) | ((s3 & k0) | ((o3 & l0) | (h3 & m0)))))))))),
  z30 = (~\[201]  & (~e19 & t2)) | ((~\[201]  & (e19 & ~t2)) | (r20 & j)),
  \[204]  = (~z50 & ~y3) | ((z50 & y3) | ~v42),
  \[7]  = (x4 & t0) | ((s4 & u0) | ((n4 & q0) | ((j4 & r0) | ((e4 & s0) | ((a4 & n0) | ((x3 & o0) | ((u3 & p0) | ((r3 & k0) | ((n3 & l0) | (g3 & m0)))))))))),
  z40 = (n40 & (~j50 & (s3 & r3))) | (n40 & (j50 & (~s3 & ~r3))),
  \[110]  = (~y50 & (~p47 & r4)) | (y50 & (~p47 & ~r4)),
  \[205]  = \[157]  | ~m2,
  \[8]  = (r5 & o0) | ((p5 & n0) | ((m5 & p0) | ((w4 & t0) | ((r4 & u0) | ((m4 & q0) | ((h4 & r0) | ((d4 & s0) | ((q3 & k0) | ((m3 & l0) | (f3 & m0)))))))))),
  z50 = ~\[146]  & ~g0,
  \[111]  = (~\[184]  & (~p47 & ~s4)) | (\[184]  & (~p47 & s4)),
  \[206]  = \[158]  | ~o4,
  \[9]  = (~\[170]  & q0) | ((k40 & m0) | ((h40 & k0) | ((~c52 & s0) | ((~e52 & o0) | ((q5 & n0) | ((n5 & p0) | ((l5 & u0) | ((v4 & t0) | ((g4 & r0) | (l3 & l0)))))))))),
  k10 = \[122] ,
  \[112]  = (~p47 & (~\[111]  & (~t4 & s4))) | ((~p47 & (t4 & ~s4)) | (\[111]  & t4)),
  k20 = (\[252]  & ~h20) | (~h20 & ~v0),
  \[113]  = (~j47 & (~p47 & (~\[112]  & t4))) | (~j47 & (~p47 & u4)),
  \[114]  = (~j47 & (~p47 & v4)) | (j47 & (~p47 & ~v4)),
  \[209]  = ~k20 & ~b,
  k40 = t3 & (s3 & (r3 & (q3 & p3))),
  \[115]  = (~\[185]  & (~p47 & ~w4)) | (\[185]  & (~p47 & w4)),
  k45 = ~\[168]  & (k4 & j4),
  \[116]  = (~p47 & (~\[115]  & (~x4 & w4))) | ((~p47 & (x4 & ~w4)) | (\[115]  & x4)),
  \[117]  = (y47 & (~p47 & (~\[116]  & x4))) | (y47 & (~p47 & y4)),
  \[118]  = (~y47 & (~p47 & ~z4)) | (y47 & (~p47 & z4)),
  \[210]  = ~l51 & ~z,
  \[211]  = o26 & ~q19,
  \[212]  = ~v50 & n44,
  \[121]  = (v49 & (~o49 & ~d5)) | e5,
  l10 = \[123] ,
  \[122]  = (g49 & (o49 & ~y48)) | (g49 & ~d5),
  \[123]  = (\[165]  & (~y48 & \[121] )) | (\[121]  & ~e5),
  \[124]  = (~\[163]  & (f50 & (~g5 & ~f5))) | ((\[163]  & (f50 & f5)) | z),
  l37 = (~\[174]  & (c52 & ~j50)) | ((~\[173]  & (c52 & j50)) | (~\[144]  & (c52 & q5))),
  \[125]  = (\[163]  & (g5 & ~z)) | ((~\[124]  & f5) | ~f50),
  l51 = (\[253]  & ~j51) | ((~j51 & u53) | ~\[241] ),
  \[126]  = (~\[170]  & (~h5 & ~z)) | ((\[170]  & (h5 & ~z)) | ~f50),
  \[128]  = (~m53 & (~k5 & ~j5)) | (m53 & (j5 & ~z)),
  \[129]  = (~m53 & (~k5 & j5)) | (\[128]  & k5),
  \[130]  = (~o49 & (~y48 & ~e52)) | ((\[195]  & ~m53) | ((~k40 & ~m53) | j51)),
  \[131]  = (~y48 & (~y47 & (~u53 & z4))) | ((~y48 & (~u53 & (~r5 & z4))) | ((~y48 & (~u53 & a0)) | ((\[195]  & ~m53) | ((~y48 & ~e52) | ~\[187] )))),
  m10 = \[124] ,
  \[132]  = (~y48 & (u53 & ~m5)) | ((~y48 & (~\[130]  & l5)) | (h40 & ~m53)),
  m16 = ~\[177]  & (y0 & (x0 & w0)),
  m19 = ~\[188]  & ~z0,
  \[133]  = ~u53,
  \[134]  = (~\[256]  & (~x53 & ~p5)) | (~\[136]  & ~\[135] ),
  \[135]  = (\[259]  & (c54 & q5)) | ((~x53 & (c54 & r5)) | (~w53 & (c54 & p5))),
  m53 = \[232]  | ~e52,
  \[136]  = (\[259]  & (c54 & r5)) | ((~x53 & (c54 & p5)) | (~w53 & (c54 & q5))),
  \[231]  = n1 | ~m1,
  \[232]  = n5 | ~m5,
  n10 = \[125] ,
  \[143]  = h22 | j,
  a6 = \[8] ,
  a7 = \[34] ,
  a8 = \[60] ,
  \[144]  = m53 | h0,
  a9 = \[86] ,
  \[239]  = ~j26 | ~g2,
  n38 = (~\[203]  & (~j50 & i3)) | ((~\[203]  & (j50 & ~i3)) | (c52 & h0)),
  n40 = (w39 & (~j50 & q3)) | (w39 & (j50 & ~q3)),
  b6 = \[9] ,
  b7 = \[35] ,
  b8 = \[61] ,
  n43 = (\[254]  & (v42 & (~z3 & ~y3))) | ((v42 & (~z50 & (z3 & y3))) | (q42 & i0)),
  \[145]  = \[21]  | g1,
  b9 = \[87] ,
  n44 = (\[243]  & ~\[183] ) | ~g4,
  n50 = ~y4 & (~x4 & (~w4 & r50)),
  c6 = \[10] ,
  c7 = \[36] ,
  c8 = \[62] ,
  \[146]  = \[121]  | c5,
  c9 = \[88] ,
  d6 = \[11] ,
  d7 = \[37] ,
  d8 = \[63] ,
  d9 = \[89] ,
  e6 = \[12] ,
  e7 = \[38] ,
  e8 = \[64] ,
  e9 = \[90] ,
  f6 = \[13] ,
  f7 = \[39] ,
  f8 = \[65] ,
  f9 = \[91] ,
  g6 = \[14] ,
  g7 = \[40] ,
  g8 = \[66] ,
  g9 = \[92] ,
  h6 = \[15] ,
  h7 = \[41] ,
  h8 = \[67] ,
  h9 = \[93] ,
  i6 = \[16] ,
  i7 = \[42] ,
  i8 = \[68] ,
  i9 = \[94] ,
  \[241]  = u53 | r4,
  j6 = \[17] ,
  j7 = \[43] ,
  j8 = \[69] ,
  j9 = \[95] ,
  k6 = \[18] ,
  k7 = \[44] ,
  k8 = \[70] ,
  k9 = \[96] ,
  \[243]  = ~i44 | ~i4,
  l6 = a,
  l7 = \[45] ,
  l8 = \[71] ,
  l9 = \[97] ,
  m6 = e1,
  m7 = \[46] ,
  m8 = \[72] ,
  m9 = \[98] ,
  n6 = \[21] ,
  n7 = \[47] ,
  n8 = \[73] ,
  n9 = \[99] ,
  o10 = \[126] ,
  o6 = \[22] ,
  o7 = \[48] ,
  o8 = \[74] ,
  o9 = \[100] ,
  \[247]  = \[181]  | ~j1,
  p6 = \[23] ,
  p7 = \[49] ,
  p8 = \[75] ,
  p9 = \[101] ,
  o26 = (\[239]  & ~\[180] ) | ~e2,
  q6 = \[24] ,
  q7 = \[50] ,
  q8 = \[76] ,
  q9 = \[102] ,
  \[249]  = \[190]  | ~e3,
  r6 = j1,
  r7 = \[51] ,
  r8 = \[77] ,
  \[155]  = l51 & ~z,
  r9 = \[103] ,
  o49 = b5 | ~a5,
  s5 = \[0] ,
  s6 = \[26] ,
  s7 = \[52] ,
  s8 = \[78] ,
  \[156]  = k20 & ~b,
  s9 = \[104] ,
  t5 = \[1] ,
  t6 = \[27] ,
  t7 = \[53] ,
  t8 = \[79] ,
  \[157]  = ~a28 | ~l2,
  t9 = \[105] ,
  u5 = \[2] ,
  u6 = \[28] ,
  u7 = \[54] ,
  u8 = \[80] ,
  \[158]  = ~b46 | ~n4,
  u9 = \[106] ,
  v5 = \[3] ,
  v6 = \[29] ,
  v7 = \[55] ,
  v8 = \[81] ,
  \[159]  = \[145]  | j18,
  v9 = \[107] ,
  w5 = \[4] ,
  w6 = \[30] ,
  w7 = \[56] ,
  w8 = \[82] ,
  w9 = \[108] ,
  x5 = \[5] ,
  x6 = \[31] ,
  x7 = \[57] ,
  x8 = \[83] ,
  x9 = \[109] ,
  y5 = \[6] ,
  y6 = \[32] ,
  y7 = \[58] ,
  y8 = \[84] ,
  y9 = \[110] ,
  z5 = \[7] ,
  z6 = \[33] ,
  z7 = \[59] ,
  z8 = \[85] ,
  z9 = \[111] ,
  \[252]  = ~i19 | (p22 | (d1 | w0)),
  \[253]  = ~n50 | (z4 | s4),
  \[254]  = q42 & ~x3,
  \[160]  = \[146]  | g49,
  \[255]  = t22,
  \[256]  = w53,
  p10 = g5,
  \[257]  = ~m1 & l1,
  p21 = ~e3 & (~d3 & (~c3 & (~b3 & (~a3 & (~z2 & y2))))),
  p22 = (n1 & ~b) | ((m1 & ~b) | h20),
  \[163]  = ~\[126]  | h5,
  p25 = (c25 & (~v19 & x1)) | ((c25 & (v19 & ~x1)) | (s24 & k)),
  \[258]  = u22 & t22,
  \[164]  = ~o1 | (k1 | ~j1),
  p36 = (\[173]  & (r36 & ~q5)) | ((\[173]  & \[144] ) | ((~r36 & ~p5) | (r36 & h3))),
  \[259]  = x53 & w53,
  \[165]  = ~o5 | (i5 | ~g5),
  p47 = (~m53 & (r5 & r4)) | ((~\[160]  & ~u53) | y48),
  \[166]  = o26 | ~f2,
  a10 = \[112] ,
  \[167]  = (j27 & j2) | l,
  a26 = (p25 & (~v19 & (z1 & y1))) | (~\[179]  & (p25 & ~z1)),
  \[168]  = n44 | ~h4,
  a28 = \[167]  & k2,
  \[169]  = (k45 & l4) | j0,
  \[260]  = z30 & e19,
  \[261]  = z30 & ~e19,
  \[262]  = n38 & j50,
  \[10]  = (~u19 & (~s16 & v0)) | (u19 & (~s16 & ~v0)),
  \[263]  = n38 & ~j50,
  \[11]  = (~\[177]  & (~s16 & ~w0)) | (\[177]  & (~s16 & w0)),
  \[12]  = (~s16 & (~\[11]  & (~x0 & w0))) | ((~s16 & (x0 & ~w0)) | (\[11]  & x0)),
  \[170]  = n44 | ~p4,
  \[13]  = (~m16 & (~s16 & (~\[12]  & x0))) | (~m16 & (~s16 & y0)),
  \[171]  = r2 | q2,
  \[14]  = (~m16 & (~s16 & z0)) | (m16 & (~s16 & ~z0)),
  q10 = \[128] ,
  \[172]  = ~r2 | ~q2,
  q19 = (b18 & t20) | ~\[181] ,
  \[15]  = (~\[178]  & (~s16 & ~a1)) | (\[178]  & (~s16 & a1)),
  \[173]  = g3 | f3,
  \[16]  = (~s16 & (~\[15]  & (~b1 & a1))) | ((~s16 & (b1 & ~a1)) | (\[15]  & b1)),
  \[174]  = ~g3 | ~f3,
  q39 = (\[263]  & k3) | (\[262]  & j3),
  \[17]  = (b17 & (~s16 & (~\[16]  & b1))) | (b17 & (~s16 & c1)),
  q42 = (~\[198]  & (~z50 & w3)) | ((~\[198]  & (z50 & ~w3)) | (~g41 & i0)),
  \[175]  = ~j50 & ~e52,
  \[18]  = (~b17 & (~s16 & ~d1)) | (b17 & (~s16 & d1)),
  \[176]  = ~e19 & ~t20,
  b10 = \[113] ,
  \[177]  = ~u19 | ~v0,
  b17 = \[178]  | (~c1 | (~b1 | ~a1)),
  b18 = (\[257]  & n1) | b,
  \[178]  = ~m16 | ~z0,
  b32 = (\[261]  & v2) | (\[260]  & u2),
  \[179]  = ~v19 | y1,
  b46 = \[169]  & m4,
  \[21]  = (y18 & (~r18 & ~h1)) | i1,
  \[22]  = (j18 & (r18 & ~b18)) | (j18 & ~h1),
  \[180]  = p1 | l,
  \[23]  = (\[164]  & (~b18 & \[21] )) | (\[21]  & ~i1),
  \[181]  = o26 | ~n2,
  \[24]  = (~q19 & (~b18 & j1)) | ((q19 & (~b18 & ~j1)) | (\[257]  & t20)),
  r10 = \[129] ,
  \[182]  = ~z50 | a4,
  r18 = f1 | ~e1,
  r20 = (~\[252]  & (\[159]  & ~v0)) | ((~h22 & ~r1) | ((~h22 & v0) | f)),
  \[183]  = p5 | j0,
  \[26]  = (~r18 & (~b18 & ~t20)) | ((\[249]  & ~h22) | ((\[191]  & ~h22) | h20)),
  \[184]  = ~y50 | ~r4,
  r36 = (\[174]  & (~q5 & ~p5)) | ((\[174]  & \[144] ) | ((\[144]  & ~h3) | (~p5 & ~h3))),
  r38 = (\[263]  & l3) | (\[262]  & ~l3),
  \[27]  = (~b18 & (~b17 & (~p22 & d1))) | ((~b18 & (~p22 & (~r1 & d1))) | ((~b18 & (~p22 & c)) | ((\[191]  & ~h22) | ((~b18 & ~t20) | ~\[186] )))),
  \[185]  = ~j47 | ~v4,
  \[28]  = (~b18 & (p22 & ~m1)) | ((~b18 & (~\[26]  & l1)) | (p21 & ~h22)),
  r50 = ~\[189]  & ~v4,
  \[186]  = b18 | ~n1,
  c10 = \[114] ,
  \[29]  = ~p22,
  \[187]  = y48 | ~n5,
  c25 = (~\[199]  & (~v19 & w1)) | (~\[199]  & (v19 & ~w1)),
  \[188]  = y0 | x0,
  \[189]  = u4 | t4,
  c52 = (~\[253]  & (~\[241]  & \[160] )) | ((~r5 & (k5 & ~j5)) | ((k5 & (~j5 & r4)) | d0)),
  c54 = (~r5 & (~q5 & ~z)) | ((~r5 & (~p5 & ~z)) | (~q5 & (~p5 & ~z))),
  \[30]  = (~\[255]  & (~u22 & ~p1)) | (~\[32]  & ~\[31] ),
  \[31]  = (\[258]  & (z22 & q1)) | ((~u22 & (z22 & r1)) | (~t22 & (z22 & p1))),
  \[32]  = (\[258]  & (z22 & r1)) | ((~u22 & (z22 & p1)) | (~t22 & (z22 & q1))),
  \[190]  = ~d3 | ~c3,
  \[33]  = (\[156]  & (~d21 & ~s1)) | ((\[156]  & (d21 & s1)) | (\[209]  & w2)),
  \[191]  = p21 | r18,
  \[34]  = (\[156]  & (~x23 & t1)) | ((\[156]  & (x23 & ~t1)) | (\[209]  & x2)),
  s10 = \[130] ,
  s16 = (~h22 & (r1 & v0)) | ((~\[159]  & ~p22) | b18),
  \[35]  = (~\[197]  & (\[156]  & ~u1)) | ((\[197]  & (\[156]  & u1)) | (\[209]  & y2)),
  \[193]  = ~c2 | ~b2,
  s24 = (~\[197]  & (~v19 & u1)) | ((~\[197]  & (v19 & ~u1)) | (~d21 & k)),
  \[36]  = (~s24 & (k20 & v1)) | ((s24 & (k20 & ~v1)) | ((~k20 & z2) | b)),
  \[194]  = ~e4 | ~d4,
  \[37]  = (~\[199]  & (k20 & ~w1)) | ((\[199]  & (k20 & w1)) | ((~k20 & a3) | b)),
  \[195]  = o49 | h40,
  \[38]  = (~c25 & (k20 & x1)) | ((c25 & (k20 & ~x1)) | ((~k20 & b3) | b)),
  d10 = \[115] ,
  \[39]  = (\[156]  & (~p25 & y1)) | ((\[156]  & (p25 & ~y1)) | (\[209]  & c3)),
  \[197]  = (~v19 & ~t1) | ((v19 & t1) | ~x23),
  d21 = (~i19 & (~q1 & (~p1 & ~h))) | ((~r1 & (~q1 & (~p1 & ~h))) | ((~m19 & (~p1 & ~h)) | ((\[188]  & ~h) | ((p22 & ~h) | ((~w0 & ~h) | (v0 & ~h)))))),
  \[198]  = (~z50 & ~v3) | ((z50 & v3) | ~v41),
  d31 = (\[261]  & w2) | (\[260]  & ~w2),
  \[199]  = (~v19 & ~v1) | ((v19 & v1) | ~s24),
  \[40]  = (~a26 & (p25 & (k20 & (~v19 & y1)))) | ((\[179]  & (~a26 & (k20 & z1))) | ((a26 & (k20 & v19)) | ((~p25 & (k20 & z1)) | ((~k20 & d3) | b)))),
  \[41]  = (~a26 & (k20 & a2)) | ((a26 & (k20 & ~a2)) | ((~k20 & e3) | b)),
  \[42]  = b | ~b2,
  \[43]  = (~c2 & b2) | ((c2 & ~b2) | b),
  \[44]  = (~\[193]  & ~d2) | ((\[193]  & d2) | b),
  t10 = \[131] ,
  \[45]  = (~\[239]  & \[211] ) | ((\[211]  & \[180] ) | ((\[211]  & e2) | ((q19 & s1) | b))),
  t20 = (\[231]  & ~b) | (l1 & ~b),
  t22 = (\[186]  & ~e) | (~l1 & ~e),
  \[46]  = (~o26 & (~q19 & ~f2)) | ((\[211]  & f2) | ((q19 & t1) | b)),
  \[47]  = (~j26 & g2) | ((j26 & ~g2) | b),
  \[48]  = (~\[166]  & (~q19 & ~h2)) | ((\[166]  & (~q19 & h2)) | ((q19 & u1) | b)),
  e10 = \[116] ,
  \[49]  = (~\[166]  & (~j27 & (~q19 & h2))) | ((~j27 & (~q19 & i2)) | ((q19 & v1) | b)),
  e19 = (~\[145]  & ~g) | (p22 & ~g),
  e29 = (\[171]  & (g29 & ~q1)) | ((\[171]  & \[143] ) | ((g29 & s2) | (s2 & ~p1))),
  e52 = (\[232]  & ~z) | (l5 & ~z),
  \[50]  = (~j27 & (~q19 & j2)) | ((j27 & (~q19 & ~j2)) | ((q19 & w1) | b)),
  \[51]  = (\[167]  & (~a28 & ~q19)) | ((~a28 & (~q19 & k2)) | ((q19 & x1) | b)),
  \[52]  = (~a28 & (~q19 & l2)) | ((a28 & (~q19 & ~l2)) | ((q19 & y1) | b)),
  \[53]  = (~\[157]  & (~q19 & ~m2)) | ((\[157]  & (~q19 & m2)) | ((q19 & z1) | b)),
  \[54]  = (~q19 & (o2 & (m2 & (l2 & (k2 & (j2 & (i2 & (h2 & f2)))))))) | (o2 & (m2 & (l2 & (k2 & (j2 & (i2 & (h2 & (f2 & b)))))))),
  u10 = \[132] ,
  u19 = (~h22 & r1) | \[159] ,
  \[55]  = (~\[205]  & (~q19 & ~o2)) | ((\[205]  & (~q19 & o2)) | ((q19 & a2) | b)),
  u22 = (\[186]  & ~d) | (m1 & ~d),
  \[56]  = (~\[247]  & ~a) | (\[247]  & p2),
  \[57]  = (~r20 & (t20 & q2)) | (r20 & (t20 & ~q2)),
  \[58]  = (~\[200]  & (t20 & ~r2)) | (\[200]  & (t20 & r2)),
  u53 = (n5 & ~z) | ((m5 & ~z) | j51),
  f10 = \[117] ,
  \[59]  = (~x29 & (t20 & s2)) | (x29 & (t20 & ~s2)),
  f50 = (~j51 & ~y48) | ~u53,
  \[60]  = (~\[201]  & (t20 & ~t2)) | ((\[201]  & (t20 & t2)) | \[176] ),
  \[61]  = (t20 & (~z2 & (~y2 & (~x2 & ~w2)))) | (e19 & ~t20),
  \[62]  = t20 & (z2 & (y2 & (x2 & w2))),
  \[63]  = (~z30 & (t20 & w2)) | (z30 & (t20 & ~w2)),
  \[64]  = (~d31 & (t20 & x2)) | (d31 & (t20 & ~x2)),
  v10 = \[133] ,
  v19 = ~\[145]  & ~i,
  \[65]  = (~h31 & (t20 & y2)) | (h31 & (t20 & ~y2)),
  \[66]  = (d31 & (~e19 & (~z2 & (y2 & x2)))) | ((d31 & (e19 & (\[64]  & (~z2 & ~y2)))) | ((e19 & (t20 & (~\[64]  & z2))) | ((~d31 & (t20 & z2)) | ((~e19 & (z2 & ~y2)) | ((\[64]  & (z2 & y2)) | \[176] ))))),
  v38 = (\[263]  & (m3 & l3)) | (\[262]  & (~m3 & ~l3)),
  \[67]  = (~b32 & (t20 & a3)) | ((b32 & (t20 & ~a3)) | \[176] ),
  v41 = (~z50 & (~g41 & u3)) | (z50 & (~g41 & ~u3)),
  v42 = (q42 & (~z50 & x3)) | (\[254]  & z50),
  v49 = \[165]  | o49,
  \[68]  = (~h32 & (t20 & b3)) | ((h32 & (t20 & ~b3)) | \[176] ),
  v50 = (y48 & e52) | ~\[170] ,
  g10 = \[118] ,
  \[69]  = (~w32 & (t20 & c3)) | (w32 & (t20 & ~c3)),
  g29 = (\[172]  & (~q1 & ~p1)) | ((\[172]  & \[143] ) | ((\[143]  & ~s2) | (~s2 & ~p1))),
  g41 = (~n50 & (~q5 & (~p5 & ~f0))) | ((~r5 & (~q5 & (~p5 & ~f0))) | ((~r50 & (~p5 & ~f0)) | ((\[241]  & ~f0) | ((\[189]  & ~f0) | (~s4 & ~f0))))),
  g49 = (~\[165]  & (v49 & ~e5)) | d5,
  \[70]  = (\[190]  & (w32 & (~e19 & c3))) | ((~i33 & (t20 & (~\[69]  & d3))) | ((\[190]  & (~e19 & d3)) | ((~\[190]  & \[69] ) | ((i33 & \[69] ) | \[176] )))),
  \[71]  = (~i33 & (t20 & e3)) | ((i33 & (t20 & ~e3)) | \[176] ),
  \[72]  = (~c52 & (e52 & f3)) | (c52 & (e52 & ~f3)),
  \[73]  = (~\[202]  & (e52 & ~g3)) | (\[202]  & (e52 & g3)),
  \[74]  = (~l37 & (e52 & h3)) | (l37 & (e52 & ~h3)),
  w10 = \[134] ,
  \[75]  = (~\[203]  & (e52 & ~i3)) | ((\[203]  & (e52 & i3)) | \[175] ),
  \[76]  = (e52 & (~o3 & (~n3 & (~m3 & ~l3)))) | (j50 & ~e52),
  w32 = (h32 & (~e19 & b3)) | (h32 & (e19 & ~b3));
endmodule

