// IWLS benchmark module "frg1" printed on Wed May 29 16:08:42 2002
module frg1(a, b, c, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, \x , y, z, a0, b0, c0, d0, e0, f0);
input
  c0,
  a,
  b,
  c,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  t,
  u,
  v,
  w,
  \x ,
  y,
  z,
  a0,
  b0;
output
  d0,
  e0,
  f0;
wire
  \[0] ,
  \[1] ,
  \[2] ;
assign
  d0 = \[0] ,
  e0 = \[1] ,
  f0 = \[2] ,
  \[0]  = (~\x  & (~w & (~u & (~t & (~s & (~p & (~o & (a & (~y & (~q & (~z & (~v & (~r & ~c))))))))))))) | ((~\x  & (~w & (~u & (~t & (~s & (~p & (~o & (~y & (~q & (~z & (~v & (~r & (e & ~c))))))))))))) | ((~m & (~u & (~t & (~s & (~p & (~o & (a & (~q & (~v & (~r & ~c)))))))))) | ((~m & (~u & (~t & (~s & (~p & (~o & (~q & (~v & (~r & (e & ~c)))))))))) | ((~\x  & (~w & (~p & (~o & (a & (~y & (~q & (~k & (~z & (~r & ~c)))))))))) | ((~\x  & (~w & (~p & (~o & (~y & (~q & (~k & (~z & (~r & (e & ~c)))))))))) | ((~\x  & (~t & (~s & (~p & (a & (~z & (~v & (~r & (~h & ~c))))))))) | ((~\x  & (~t & (~s & (~p & (~z & (~v & (~r & (~h & (e & ~c))))))))) | ((~i & (~\x  & (~w & (~t & (~s & (~p & (~o & (a & ~c)))))))) | ((~i & (~\x  & (~w & (~t & (~s & (~p & (~o & (e & ~c)))))))) | ((~m & (~t & (~s & (~p & (a & (~v & (~r & (~h & ~c)))))))) | ((~m & (~t & (~s & (~p & (~v & (~r & (~h & (e & ~c)))))))) | ((~u & (a & (~y & (~q & (~z & (~v & (~r & (~j & ~c)))))))) | ((~u & (~y & (~q & (~z & (~v & (~r & (~j & (e & ~c)))))))) | ((~i & (~m & (~t & (~s & (~p & (~o & (a & ~c))))))) | ((~i & (~m & (~t & (~s & (~p & (~o & (e & ~c))))))) | ((~i & (~m & (~t & (~s & (~p & (a & (~h & ~c))))))) | ((~i & (~m & (~t & (~s & (~p & (~h & (e & ~c))))))) | ((~i & (~\x  & (~w & (~p & (~o & (a & (~k & ~c))))))) | ((~i & (~\x  & (~w & (~p & (~o & (~k & (e & ~c))))))) | ((~i & (~\x  & (~t & (~s & (~p & (a & (~h & ~c))))))) | ((~i & (~\x  & (~t & (~s & (~p & (~h & (e & ~c))))))) | ((~m & (~u & (a & (~q & (~v & (~r & (~j & ~c))))))) | ((~m & (~u & (~q & (~v & (~r & (~j & (e & ~c))))))) | ((~m & (~p & (~o & (a & (~q & (~k & (~r & ~c))))))) | ((~m & (~p & (~o & (~q & (~k & (~r & (e & ~c))))))) | ((~\x  & (~p & (a & (~k & (~z & (~r & (~h & ~c))))))) | ((~\x  & (~p & (~k & (~z & (~r & (~h & (e & ~c))))))) | ((~w & (~u & (~o & (a & (~y & (~q & (~g & ~c))))))) | ((~w & (~u & (~o & (~y & (~q & (~g & (e & ~c))))))) | ((~w & (~o & (a & (~y & (~q & (~k & (~g & ~c))))))) | ((~w & (~o & (~y & (~q & (~k & (~g & (e & ~c))))))) | ((a & (~y & (~q & (~k & (~z & (~r & (~j & ~c))))))) | ((~y & (~q & (~k & (~z & (~r & (~j & (e & ~c))))))) | ((~n & (~\x  & (~w & (a & (~y & (~z & ~c)))))) | ((~n & (~\x  & (~w & (~y & (~z & (e & ~c)))))) | ((~l & (~u & (~t & (~s & (a & (~v & ~c)))))) | ((~l & (~u & (~t & (~s & (~v & (e & ~c)))))) | ((~l & (~t & (~s & (a & (~v & (~h & ~c)))))) | ((~l & (~t & (~s & (~v & (~h & (e & ~c)))))) | ((~i & (~m & (~p & (~o & (a & (~k & ~c)))))) | ((~i & (~m & (~p & (~o & (~k & (e & ~c)))))) | ((~i & (~m & (~p & (a & (~k & (~h & ~c)))))) | ((~i & (~m & (~p & (~k & (~h & (e & ~c)))))) | ((~i & (~\x  & (~p & (a & (~k & (~h & ~c)))))) | ((~i & (~\x  & (~p & (~k & (~h & (e & ~c)))))) | ((~m & (~u & (~o & (a & (~q & (~g & ~c)))))) | ((~m & (~u & (~o & (~q & (~g & (e & ~c)))))) | ((~m & (~u & (a & (~q & (~g & (~j & ~c)))))) | ((~m & (~u & (~q & (~g & (~j & (e & ~c)))))) | ((~m & (~p & (a & (~k & (~r & (~h & ~c)))))) | ((~m & (~p & (~k & (~r & (~h & (e & ~c)))))) | ((~m & (~o & (a & (~q & (~k & (~g & ~c)))))) | ((~m & (~o & (~q & (~k & (~g & (e & ~c)))))) | ((~m & (a & (~q & (~k & (~g & (~j & ~c)))))) | ((~m & (a & (~q & (~k & (~r & (~j & ~c)))))) | ((~m & (a & (~k & (~r & (~j & (~h & ~c)))))) | ((~m & (a & (~v & (~r & (~j & (~h & ~c)))))) | ((~m & (~q & (~k & (~g & (~j & (e & ~c)))))) | ((~m & (~q & (~k & (~r & (~j & (e & ~c)))))) | ((~m & (~k & (~r & (~j & (~h & (e & ~c)))))) | ((~m & (~v & (~r & (~j & (~h & (e & ~c)))))) | ((~u & (a & (~y & (~q & (~g & (~j & ~c)))))) | ((~u & (~y & (~q & (~g & (~j & (e & ~c)))))) | ((a & (~y & (~q & (~k & (~g & (~j & ~c)))))) | ((a & (~k & (~z & (~r & (~j & (~h & ~c)))))) | ((a & (~z & (~v & (~r & (~j & (~h & ~c)))))) | ((~y & (~q & (~k & (~g & (~j & (e & ~c)))))) | ((~k & (~z & (~r & (~j & (~h & (e & ~c)))))) | ((~z & (~v & (~r & (~j & (~h & (e & ~c)))))) | ((~n & (~i & (~\x  & (~w & (a & ~c))))) | ((~n & (~i & (~\x  & (~w & (e & ~c))))) | ((~n & (~i & (~\x  & (a & (~h & ~c))))) | ((~n & (~i & (~\x  & (~h & (e & ~c))))) | ((~n & (~i & (~w & (a & (~g & ~c))))) | ((~n & (~i & (~w & (~g & (e & ~c))))) | ((~n & (~\x  & (a & (~z & (~h & ~c))))) | ((~n & (~\x  & (~z & (~h & (e & ~c))))) | ((~n & (~w & (a & (~y & (~g & ~c))))) | ((~n & (~w & (~y & (~g & (e & ~c))))) | ((~n & (a & (~y & (~g & (~j & ~c))))) | ((~n & (a & (~y & (~z & (~j & ~c))))) | ((~n & (a & (~z & (~j & (~h & ~c))))) | ((~n & (~y & (~g & (~j & (e & ~c))))) | ((~n & (~y & (~z & (~j & (e & ~c))))) | ((~n & (~z & (~j & (~h & (e & ~c))))) | ((~l & (~i & (~t & (~s & (a & ~c))))) | ((~l & (~i & (~t & (~s & (e & ~c))))) | ((~l & (~u & (a & (~v & (~j & ~c))))) | ((~l & (~u & (~v & (~j & (e & ~c))))) | ((~l & (a & (~v & (~j & (~h & ~c))))) | ((~l & (~v & (~j & (~h & (e & ~c))))) | ((~i & (~m & (~o & (a & (~g & ~c))))) | ((~i & (~m & (~o & (~g & (e & ~c))))) | ((~i & (~w & (~o & (a & (~g & ~c))))) | ((~i & (~w & (~o & (~g & (e & ~c))))) | ((~l & (~i & (a & (~g & ~c)))) | ((~l & (~i & (~g & (e & ~c)))) | ((~l & (~u & (a & (~g & ~c)))) | ((~l & (~u & (~g & (e & ~c)))) | ((~c0 & (~a & (~e & ~c))) | ((~n & (~l & (a & ~c))) | ((~n & (~l & (e & ~c))) | ((~n & (~m & (a & ~c))) | ((~n & (~m & (e & ~c))) | ((~l & (a & (~k & ~c))) | ((~l & (~k & (e & ~c))) | ((~i & (a & (~j & ~c))) | ((~i & (~j & (e & ~c))) | ((a & (~g & (~h & ~c))) | ((~g & (~h & (e & ~c))) | (~b & c))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))),
  \[1]  = (e & f) | ((~a0 & f) | (c | a)),
  \[2]  = (c & ~e) | ((~b0 & ~e) | (~e & a));
endmodule

