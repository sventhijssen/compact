// IWLS benchmark module "x1" printed on Wed May 29 16:25:48 2002
module x1(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2, b2, c2, d2, e2, f2, g2, h2, i2);
input
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  t,
  u,
  v,
  w,
  y,
  z,
  a0,
  b0,
  c0,
  d0,
  e0,
  f0,
  g0,
  h0,
  i0,
  j0,
  k0,
  l0,
  m0,
  n0,
  o0,
  p0,
  q0,
  r0,
  s0,
  t0,
  u0,
  v0,
  w0,
  x0,
  y0,
  z0;
output
  a1,
  a2,
  b1,
  b2,
  c1,
  c2,
  d1,
  d2,
  e1,
  e2,
  f1,
  f2,
  g1,
  g2,
  h1,
  h2,
  i1,
  i2,
  j1,
  k1,
  l1,
  m1,
  n1,
  o1,
  p1,
  q1,
  r1,
  s1,
  t1,
  u1,
  v1,
  w1,
  x1,
  y1,
  z1;
wire
  \[5] ,
  \[6] ,
  \[46] ,
  \[7] ,
  \[47] ,
  \[48] ,
  \[75] ,
  \[21] ,
  \[76] ,
  \[22] ,
  \[77] ,
  \[23] ,
  \[78] ,
  \[24] ,
  \[25] ,
  \[50] ,
  \[26] ,
  \[51] ,
  \[27] ,
  \[29] ,
  \[54] ,
  \[55] ,
  \[56] ,
  \[58] ,
  \[30] ,
  \[31] ,
  \[32] ,
  \[33] ,
  \[34] ,
  \[35] ,
  \[36] ,
  \[61] ,
  \[37] ,
  \[38] ,
  \[39] ,
  \[10] ,
  \[65] ,
  \[11] ,
  \[66] ,
  \[12] ,
  \[67] ,
  \[13] ,
  \[14] ,
  \[0] ,
  \[40] ,
  \[1] ,
  \[41] ,
  \[17] ,
  \[2] ,
  \[42] ,
  \[18] ,
  \[3] ,
  \[4] ;
assign
  \[5]  = (\[67]  & (~\[35]  & e0)) | ((q0 & (~q & ~i)) | ((q0 & (~q & ~g)) | ((q0 & (~o & ~i)) | (q0 & (~o & ~g))))),
  \[6]  = (\[42]  & (\[39]  & (\[36]  & (p0 & (~i & (~h & ~a)))))) | ((\[67]  & (\[50]  & (~\[42]  & (\[39]  & (\[36]  & p0))))) | ((\[51]  & (\[42]  & (~\[35]  & d0))) | ((\[51]  & (~\[37]  & (~\[35]  & d0))) | ((v0 & o0) | (d0 & v))))),
  \[46]  = (\[36]  & (q0 & (~v & g))) | ((\[36]  & (p0 & g)) | (p0 & v)),
  \[7]  = \[54]  & (~\[41]  & (h & ~a)),
  \[47]  = ~\[41]  & ~\[38] ,
  \[48]  = ~l | ~b,
  \[75]  = \[47]  & o,
  \[21]  = (~\[38]  & (g0 & (~j & ~f))) | ((\[65]  & (~\[40]  & ~r)) | ((~\[40]  & (~\[38]  & g0)) | (\[77]  & n))),
  \[76]  = g0 & j,
  \[22]  = (~\[39]  & k0) | (~\[39]  & a0),
  \[77]  = \[66]  & \[65] ,
  \[23]  = ~\[24] ,
  \[78]  = ~v & ~p,
  \[24]  = (~\[61]  & (~\[26]  & ~g0)) | (~\[61]  & j),
  \[25]  = c0 | d0,
  \[50]  = ~d | ~c,
  \[26]  = r0 | f0,
  \[51]  = v | ~m,
  \[27]  = (\[78]  & (\[75]  & p0)) | ((\[78]  & (\[75]  & e0)) | ((\[75]  & (~\[42]  & p0)) | (\[75]  & (~\[42]  & e0)))),
  \[29]  = (\[46]  & (i & ~a)) | (\[61]  | (i0 | y)),
  \[54]  = (e0 & ~o) | ((d0 & ~d) | (s0 | p0)),
  a1 = \[0] ,
  a2 = \[26] ,
  \[55]  = d0 & d,
  b1 = \[1] ,
  b2 = \[27] ,
  \[56]  = ~t | ~a,
  c1 = \[2] ,
  c2 = h0,
  d1 = \[3] ,
  d2 = \[29] ,
  \[58]  = \[48]  | n,
  e1 = \[4] ,
  e2 = \[30] ,
  f1 = \[5] ,
  f2 = \[31] ,
  g1 = \[6] ,
  \[30]  = ~\[29] ,
  g2 = \[32] ,
  h1 = \[7] ,
  \[31]  = ~\[32] ,
  h2 = \[33] ,
  i1 = m0,
  \[32]  = (~z0 & (a0 & ~r)) | ((~z0 & (a0 & m)) | ((~z0 & (a0 & j)) | ((\[54]  & h) | ((\[48]  & a0) | (\[26]  | (\[18]  | (x0 | m0))))))),
  i2 = \[34] ,
  j1 = n0,
  \[33]  = ~\[34] ,
  k1 = \[10] ,
  \[34]  = (~\[58]  & (\[40]  & (~\[38]  & a0))) | ((\[77]  & ~\[58] ) | ((\[76]  & c) | ((i0 & i) | ((d0 & ~h) | (\[61]  | (\[55]  | (c0 | (b0 | y)))))))),
  l1 = \[11] ,
  \[35]  = ~p | ~o,
  m1 = \[12] ,
  \[36]  = \[35]  | ~q,
  \[61]  = h0 | z,
  n1 = \[13] ,
  \[37]  = u | e,
  o1 = \[14] ,
  \[38]  = m | a,
  p1 = y,
  \[39]  = ~s | ~r,
  q1 = z,
  \[10]  = (\[55]  & (w & ~v)) | ((g0 & (~j & a)) | ((~\[56]  & i0) | ((~\[51]  & \[25] ) | ((~\[51]  & p0) | ((~\[39]  & p0) | ((~\[39]  & l0) | ((\[38]  & s0) | ((\[38]  & q0) | ((\[38]  & k0) | ((\[38]  & h0) | ((\[38]  & e0) | ((~\[2]  & b0) | ((r0 & b) | ((p0 & a) | ((j0 & a) | ((g0 & m) | ((d0 & a) | (a0 & a)))))))))))))))))),
  \[65]  = ~\[38]  & k0,
  r1 = \[17] ,
  \[11]  = (\[78]  & (\[55]  & (\[37]  & (o & ~a)))) | ((\[78]  & (\[37]  & (e0 & (o & ~a)))) | ((~\[42]  & (\[37]  & (~\[35]  & (d0 & ~a)))) | ((\[55]  & (~\[42]  & (\[37]  & ~a))) | ((~\[42]  & (\[37]  & (e0 & ~a))) | ((\[37]  & (e0 & h)) | ((\[37]  & (d0 & h)) | ((a0 & (k & b)) | ((\[41]  & h0) | ((~\[36]  & q0) | ((~\[36]  & p0) | (f0 & b))))))))))),
  \[66]  = v & ~j,
  s1 = \[18] ,
  \[12]  = (\[78]  & (\[75]  & \[55] )) | (h0 & j),
  \[67]  = ~\[38]  & ~h,
  t1 = x0,
  \[13]  = (\[47]  & (~\[35]  & (q0 & (~q & ~g)))) | ((\[66]  & (g0 & (f & ~a))) | ((~\[50]  & (\[47]  & (~\[42]  & p0))) | ((\[76]  & (\[67]  & ~c)) | ((\[75]  & (e0 & ~p)) | ((\[47]  & (w0 & o0)) | ((\[47]  & (s0 & ~h)) | (\[47]  & (h0 & ~j)))))))),
  u1 = y0,
  \[14]  = (i0 & (i & (~h & ~a))) | (\[46]  & (i & ~a)),
  v1 = \[21] ,
  \[0]  = (~\[40]  & (a0 & ~r)) | ((\[58]  & a0) | ((\[26]  & ~b) | (a0 & m))),
  w1 = \[22] ,
  \[40]  = v | j,
  \[1]  = (~\[58]  & (\[40]  & (~\[38]  & (a0 & ~k)))) | ((\[77]  & (~n & b)) | ((\[76]  & (~w & c)) | (t0 & o0))),
  x1 = \[23] ,
  \[41]  = \[37]  | w,
  \[17]  = (~\[48]  & (~\[40]  & (\[39]  & (~\[38]  & (a0 & (r & ~k)))))) | ((\[65]  & (~\[40]  & (\[39]  & (r & b)))) | ((\[56]  & (i0 & (~i & ~h))) | (j0 & ~a))),
  \[2]  = \[51]  & b0,
  y1 = \[24] ,
  \[42]  = v | g,
  \[18]  = i0 & (t & h),
  \[3]  = (\[67]  & (\[35]  & (d0 & (~v & ~d)))) | (\[51]  & c0),
  z1 = \[25] ,
  \[4]  = (\[55]  & (\[37]  & (~o & (~m & g)))) | ((\[55]  & (~\[41]  & (~o & ~m))) | ((\[67]  & (e0 & ~o)) | (u0 & o0)));
endmodule

