// IWLS benchmark module "f51m" printed on Wed May 29 16:08:42 2002
module f51m(\1 , \2 , \3 , \4 , \5 , \6 , \7 , \8 , \44 , \45 , \46 , \47 , \48 , \49 , \50 , \51 );
input
  \1 ,
  \2 ,
  \3 ,
  \4 ,
  \5 ,
  \6 ,
  \7 ,
  \8 ;
output
  \44 ,
  \45 ,
  \46 ,
  \47 ,
  \48 ,
  \49 ,
  \50 ,
  \51 ;
wire
  \[7] ,
  \[8] ,
  \[1] ,
  \[2] ,
  \[3] ,
  \[4] ,
  \[5] ,
  \[6] ;
assign
  \[7]  = (~\8  & \7 ) | (\8  & ~\7 ),
  \[8]  = ~\8 ,
  \[1]  = (~\8  & (~\6  & (~\5  & (\3  & (~\2  & ~\1 ))))) | ((\8  & (\7  & (\6  & (\3  & (\2  & \1 ))))) | ((\8  & (\6  & (\5  & (~\3  & (\2  & ~\1 ))))) | ((~\7  & (~\6  & (~\5  & (\3  & (~\2  & ~\1 ))))) | ((\7  & (\6  & (\5  & (~\3  & (\2  & ~\1 ))))) | ((~\8  & (~\7  & (~\4  & (~\3  & \1 )))) | ((~\8  & (~\5  & (~\4  & (\3  & ~\1 )))) | ((\8  & (\7  & (\4  & (\3  & \1 )))) | ((~\7  & (~\6  & (~\3  & (~\2  & \1 )))) | ((~\7  & (~\5  & (~\4  & (\3  & ~\1 )))) | ((\7  & (\5  & (\4  & (~\3  & ~\1 )))) | ((~\6  & (~\5  & (~\4  & (\3  & ~\1 )))) | ((\6  & (\5  & (\4  & (~\3  & ~\1 )))) | ((~\6  & (~\4  & (~\3  & \1 ))) | ((\6  & (\4  & (\3  & \1 ))) | ((~\5  & (~\4  & (~\3  & \1 ))) | ((~\5  & (~\3  & (~\2  & \1 ))) | ((\5  & (\4  & (\3  & \1 ))) | ((\5  & (\3  & (\2  & \1 ))) | ((~\4  & (~\3  & (~\2  & \1 ))) | ((~\4  & (\3  & (~\2  & ~\1 ))) | ((\4  & (~\3  & (\2  & ~\1 ))) | (\4  & (\3  & (\2  & \1 )))))))))))))))))))))))),
  \[2]  = (\8  & (\7  & (~\6  & (~\5  & (\3  & \2 ))))) | ((\8  & (\7  & (\6  & (~\4  & (\3  & ~\2 ))))) | ((~\8  & (~\7  & (~\4  & (~\3  & \2 )))) | ((~\8  & (~\6  & (~\5  & (\4  & ~\2 )))) | ((\8  & (\6  & (\5  & (~\4  & ~\2 )))) | ((~\7  & (~\6  & (~\5  & (\4  & ~\2 )))) | ((~\7  & (~\6  & (\4  & (~\3  & ~\2 )))) | ((\7  & (\6  & (\5  & (~\4  & ~\2 )))) | ((~\8  & (~\5  & (~\4  & \2 ))) | ((~\7  & (~\5  & (~\4  & \2 ))) | ((\7  & (\5  & (\4  & \2 ))) | ((~\6  & (~\4  & (~\3  & \2 ))) | ((\6  & (\5  & (\4  & \2 ))) | ((\6  & (\4  & (\3  & \2 ))) | ((~\5  & (~\4  & (~\3  & \2 ))) | ((~\5  & (\4  & (~\3  & ~\2 ))) | ((\5  & (~\4  & (\3  & ~\2 ))) | (\5  & (\4  & (\3  & \2 ))))))))))))))))))),
  \[3]  = (~\8  & (~\7  & (\5  & (~\4  & ~\3 )))) | ((\8  & (~\7  & (\6  & (~\4  & \3 )))) | ((\8  & (\7  & (\6  & (~\5  & ~\3 )))) | ((\8  & (\7  & (~\5  & (\4  & ~\3 )))) | ((~\8  & (~\6  & (~\5  & \3 ))) | ((~\8  & (~\5  & (~\4  & \3 ))) | ((~\7  & (~\6  & (~\5  & \3 ))) | ((~\7  & (~\6  & (\5  & ~\3 ))) | ((\7  & (\6  & (\5  & \3 ))) | ((\7  & (\5  & (\4  & \3 ))) | ((~\6  & (~\5  & (~\4  & \3 ))) | ((~\6  & (\5  & (~\4  & ~\3 ))) | ((\6  & (~\5  & (\4  & ~\3 ))) | (\6  & (\5  & (\4  & \3 ))))))))))))))),
  \[4]  = (~\8  & (~\7  & (\6  & ~\4 ))) | ((~\8  & (~\6  & (~\5  & \4 ))) | ((~\8  & (\6  & (~\5  & ~\4 ))) | ((\8  & (~\7  & (\5  & \4 ))) | ((\8  & (\7  & (~\6  & ~\4 ))) | ((\8  & (\7  & (\6  & \4 ))) | ((~\7  & (\6  & (~\5  & ~\4 ))) | ((\7  & (~\6  & (\5  & ~\4 ))) | ((\7  & (\6  & (\5  & \4 ))) | (~\7  & (~\6  & \4 )))))))))),
  \44  = \[1] ,
  \45  = \[2] ,
  \46  = \[3] ,
  \47  = \[4] ,
  \48  = \[5] ,
  \[5]  = (\8  & (~\7  & (\6  & ~\5 ))) | ((~\8  & (~\7  & \5 )) | ((~\8  & (\7  & ~\5 )) | ((\8  & (\7  & \5 )) | (~\7  & (~\6  & \5 ))))),
  \49  = \[6] ,
  \50  = \[7] ,
  \51  = \[8] ,
  \[6]  = (\8  & (~\7  & ~\6 )) | ((~\8  & \6 ) | (\7  & \6 ));
endmodule

