module foobar(z7, a8, b8, c8, d8, e8, f8, g8, h8, i8, j8, k8, l8, m8, n8, o8, p8, q8, r8, s8, t8, u8, v8, w8, x8, y8, z8, a9, b9, c9, d9, e9, f9, g9, h9, i9, j9, k9, l9, m9, n9, o9, p9, q9, r9, s9, t9, u9, v9, w9, x9, y9, z9, a10, b10, c10, d10, e10, f10, g10, h10, i10, j10, k10, l10, m10, n10, o10, p10, q10, r10, s10, t10, u10, v10, w10, x10, y10, z10, a11, b11, c11, d11, e11, f11, g11, h11, i11, j11, k11, l11, m11, n11, o11, p11, q11, r11, s11, t11, u11, v11, w11, x11, y11, z11, a12, b12, c12, d12, e12, f12, g12, h12, i12, j12, k12, l12, m12, n12, o12, p12, q12, r12, s12, t12, u12, v12, w12, x12, y12, z12, a13, b13, c13, d13, e13, f13, g13, h13, i13, a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2, b2, c2, d2, e2, f2, g2, h2, i2, j2, k2, l2, m2, n2, o2, p2, q2, r2, s2, t2, u2, v2, w2, x2, y2, z2, a3, b3, c3, d3, e3, f3, g3, h3, i3, j3, k3, l3, m3, n3, o3, p3, q3, r3, s3, t3, u3, v3, w3, x3, y3, z3, a4, b4, c4, d4, e4, f4, g4, h4, i4, j4, k4, l4, m4, n4, o4, p4, q4, r4, s4, t4, u4, v4, w4, x4, y4, z4, a5, b5, c5, d5, e5, f5, g5, h5, i5, j5, k5, l5, m5, n5, o5, p5, q5, r5, s5, t5, u5, v5, w5, x5, y5, z5, a6, b6, c6, d6, e6, f6, g6, h6, i6, j6, k6, l6, m6, n6, o6, p6, q6, r6, s6, t6, u6, v6, w6, x6, y6, z6, a7, b7, c7, d7, e7, f7, g7, h7, i7, j7, k7, l7, m7, n7, o7, p7, q7, r7, s7, t7, u7, v7, w7, x7, y7);
input a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2, b2, c2, d2, e2, f2, g2, h2, i2, j2, k2, l2, m2, n2, o2, p2, q2, r2, s2, t2, u2, v2, w2, x2, y2, z2, a3, b3, c3, d3, e3, f3, g3, h3, i3, j3, k3, l3, m3, n3, o3, p3, q3, r3, s3, t3, u3, v3, w3, x3, y3, z3, a4, b4, c4, d4, e4, f4, g4, h4, i4, j4, k4, l4, m4, n4, o4, p4, q4, r4, s4, t4, u4, v4, w4, x4, y4, z4, a5, b5, c5, d5, e5, f5, g5, h5, i5, j5, k5, l5, m5, n5, o5, p5, q5, r5, s5, t5, u5, v5, w5, x5, y5, z5, a6, b6, c6, d6, e6, f6, g6, h6, i6, j6, k6, l6, m6, n6, o6, p6, q6, r6, s6, t6, u6, v6, w6, x6, y6, z6, a7, b7, c7, d7, e7, f7, g7, h7, i7, j7, k7, l7, m7, n7, o7, p7, q7, r7, s7, t7, u7, v7, w7, x7, y7;
output z7, a8, b8, c8, d8, e8, f8, g8, h8, i8, j8, k8, l8, m8, n8, o8, p8, q8, r8, s8, t8, u8, v8, w8, x8, y8, z8, a9, b9, c9, d9, e9, f9, g9, h9, i9, j9, k9, l9, m9, n9, o9, p9, q9, r9, s9, t9, u9, v9, w9, x9, y9, z9, a10, b10, c10, d10, e10, f10, g10, h10, i10, j10, k10, l10, m10, n10, o10, p10, q10, r10, s10, t10, u10, v10, w10, x10, y10, z10, a11, b11, c11, d11, e11, f11, g11, h11, i11, j11, k11, l11, m11, n11, o11, p11, q11, r11, s11, t11, u11, v11, w11, x11, y11, z11, a12, b12, c12, d12, e12, f12, g12, h12, i12, j12, k12, l12, m12, n12, o12, p12, q12, r12, s12, t12, u12, v12, w12, x12, y12, z12, a13, b13, c13, d13, e13, f13, g13, h13, i13;
not(f11, f0);
not(g11, b3);
not(h11, l1);
not(i11, x1);
not(j11, a1);
not(k11, r2);
not(l11, q0);
not(m11, h2);
not(n11, p15);
not(o11, j17);
and(q11, v1, p11);
not(r11, i17);
not(t_0, i17);
not(t_1, m6);
or(s11, t_0, t_1);
not(t11, v17);
not(v11, u11);
not(x11, f26);
not(y11, g26);
not(z11, e26);
not(a12, o26);
not(b12, n26);
not(c12, m26);
or(d12, s27, q16);
not(e12, k31);
not(f12, g30);
or(r12, t27, g33);
not(t_2, y40);
not(t_3, v40);
or(u12, t_2, t_3);
not(w12, i46);
not(x12, k46);
not(z12, y12);
or(a13, u27, r54);
not(g13, x57);
not(i13, h13);
not(p14, y7);
not(q14, x7);
not(r14, w7);
not(s14, v7);
not(t14, u7);
not(u14, t7);
not(v14, s7);
not(w14, r7);
not(x14, q7);
not(y14, p7);
buf(z14, n7);
buf(a15, n7);
buf(b15, m7);
buf(c15, m7);
not(d15, l7);
buf(e15, l7);
not(f15, k7);
buf(g15, k7);
not(h15, j7);
buf(i15, j7);
not(j15, i7);
buf(k15, i7);
not(l15, h7);
buf(m15, h7);
not(n15, g7);
buf(o15, g7);
and(p15, j7, i7, h7, g7);
not(q15, f7);
buf(r15, f7);
not(s15, d7);
buf(t15, d7);
not(u15, c7);
buf(v15, c7);
not(w15, b7);
buf(x15, b7);
not(y15, a7);
buf(z15, a7);
not(a16, z6);
buf(b16, z6);
not(c16, y6);
buf(d16, y6);
not(e16, x6);
buf(f16, x6);
not(g16, w6);
buf(h16, w6);
not(i16, v6);
buf(j16, v6);
not(k16, u6);
not(l16, t6);
buf(m16, t6);
not(n16, s6);
buf(o16, s6);
not(p16, q6);
not(q16, p6);
buf(r16, o6);
buf(s16, n6);
buf(t16, n6);
not(u16, l6);
buf(v16, k6);
buf(w16, k6);
buf(p11, i6);
and(y16, r2, q0, h2, a1);
and(z16, b3, l1, x1, f0);
buf(a17, c0);
buf(b17, w);
buf(c17, w);
buf(d17, l);
buf(e17, l);
and(f17, i, q6);
buf(g17, h);
buf(h17, h);
and(i17, g, o6);
and(j17, b, k, o6);
and(k17, a, c);
not(t_4, p14);
not(t_5, r15);
or(l17, t_4, t_5);
not(t_6, q14);
not(t_7, j16);
or(m17, t_6, t_7);
not(t_8, s14);
not(t_9, w7);
or(n17, t_8, t_9);
not(t_10, r14);
not(t_11, v7);
or(o17, t_10, t_11);
not(t_12, u14);
not(t_13, u7);
or(p17, t_12, t_13);
not(t_14, t14);
not(t_15, t7);
or(q17, t_14, t_15);
not(t_16, w14);
not(t_17, s7);
or(r17, t_16, t_17);
not(t_18, v14);
not(t_19, r7);
or(s17, t_18, t_19);
not(t_20, y14);
not(t_21, q7);
or(t17, t_20, t_21);
not(t_22, x14);
not(t_23, p7);
or(u17, t_22, t_23);
and(v17, o7, i17);
not(w17, z14);
and(x17, c15, a15);
not(y17, a15);
not(z17, b15);
not(a18, c15);
not(b18, e15);
not(c18, g15);
buf(d18, h15);
not(e18, i15);
buf(f18, j15);
not(g18, k15);
buf(h18, l15);
not(i18, m15);
buf(j18, n15);
not(k18, o15);
buf(l18, q15);
not(m18, r15);
buf(n18, s15);
not(o18, t15);
buf(p18, u15);
not(q18, v15);
buf(r18, w15);
not(s18, x15);
buf(t18, y15);
not(u18, z15);
buf(v18, a16);
not(w18, b16);
buf(x18, c16);
not(y18, d16);
buf(z18, e16);
not(a19, f16);
buf(b19, g16);
not(c19, h16);
buf(d19, i16);
not(e19, j16);
buf(f19, l16);
not(g19, m16);
buf(h19, n16);
not(i19, o16);
not(j19, s16);
not(k19, t16);
not(l19, v16);
not(m19, w16);
and(n19, p2, b15, z14);
and(o19, o2, b15, z14);
and(p19, n2, b15, z14);
and(q19, m2, b15, z14);
and(r19, l2, c15, a15);
and(s19, k2, c15, a15);
and(t19, j2, c15, a15);
and(u19, i2, c15, a15);
and(v19, g2, b15, z14);
and(w19, j1, w16, t16);
and(x19, i1, w16, t16);
and(y19, h1, w16, t16);
and(z19, g1, w16, t16);
and(a20, f1, v16, s16);
and(b20, e1, v16, s16);
and(c20, d1, v16, s16);
and(d20, c1, v16, s16);
and(e20, b1, v16, s16);
and(f20, z0, w16, t16);
and(u11, y16, z16);
not(h20, y16);
not(i20, z16);
not(j20, a17);
not(k20, b17);
not(l20, c17);
not(m20, d17);
not(n20, e17);
and(o20, i, p16);
buf(p20, g17);
buf(q20, g17);
buf(r20, h17);
buf(s20, h17);
not(t20, k17);
not(t_24, m18);
not(t_25, y7);
or(u20, t_24, t_25);
not(t_26, e19);
not(t_27, x7);
or(v20, t_26, t_27);
not(t_28, o17);
not(t_29, n17);
or(w20, t_28, t_29);
not(t_30, q17);
not(t_31, p17);
or(x20, t_30, t_31);
not(t_32, s17);
not(t_33, r17);
or(y20, t_32, t_33);
not(t_34, u17);
not(t_35, t17);
or(z20, t_34, t_35);
and(a21, o7, i20);
and(b21, a18, a15);
and(c21, a18, y17);
and(d21, c15, y17);
not(t_36, c18);
not(t_37, e15);
or(e21, t_36, t_37);
not(t_38, b18);
not(t_39, g15);
or(f21, t_38, t_39);
not(g21, d18);
not(t_40, g18);
not(t_41, i15);
or(h21, t_40, t_41);
not(i21, f18);
not(t_42, e18);
not(t_43, k15);
or(j21, t_42, t_43);
not(k21, h18);
not(t_44, k18);
not(t_45, m15);
or(l21, t_44, t_45);
not(m21, j18);
not(t_46, i18);
not(t_47, o15);
or(n21, t_46, t_47);
not(o21, l18);
not(p21, n18);
not(t_48, q18);
not(t_49, t15);
or(q21, t_48, t_49);
not(r21, p18);
not(t_50, o18);
not(t_51, v15);
or(s21, t_50, t_51);
not(t21, r18);
not(t_52, u18);
not(t_53, x15);
or(u21, t_52, t_53);
not(v21, t18);
not(t_54, s18);
not(t_55, z15);
or(w21, t_54, t_55);
not(x21, v18);
not(t_56, y18);
not(t_57, b16);
or(y21, t_56, t_57);
not(z21, x18);
not(t_58, w18);
not(t_59, d16);
or(a22, t_58, t_59);
not(b22, z18);
not(t_60, c19);
not(t_61, f16);
or(c22, t_60, t_61);
not(d22, b19);
not(t_62, a19);
not(t_63, h16);
or(e22, t_62, t_63);
not(f22, d19);
not(g22, f19);
not(t_64, i19);
not(t_65, m16);
or(h22, t_64, t_65);
not(i22, h19);
not(t_66, g19);
not(t_67, o16);
or(j22, t_66, t_67);
and(k22, l19, s16);
and(l22, m6, h20);
and(m22, j3, z17, w17);
and(n22, i3, z17, w17);
and(o22, h3, z17, w17);
and(p22, g3, z17, w17);
and(q22, f3, a18, y17);
and(r22, e3, a18, y17);
and(s22, d3, a18, y17);
and(t22, c3, a18, y17);
and(u22, a3, z17, w17);
and(v22, z2, z17, z14);
and(w22, y2, z17, z14);
and(x22, x2, z17, z14);
and(y22, w2, z17, z14);
and(z22, v2, a18, a15);
and(a23, u2, a18, a15);
and(b23, t2, a18, a15);
and(c23, s2, a18, a15);
and(d23, q2, z17, z14);
and(e23, f2, b15, w17);
and(f23, e2, b15, w17);
and(g23, d2, b15, w17);
and(h23, c2, b15, w17);
and(i23, b2, c15, y17);
and(j23, a2, c15, y17);
and(k23, z1, c15, y17);
and(l23, y1, c15, y17);
and(m23, w1, b15, w17);
and(n23, u1, m19, k19);
and(o23, t1, m19, k19);
and(p23, s1, m19, k19);
and(q23, r1, m19, k19);
and(r23, q1, l19, j19);
and(s23, p1, l19, j19);
and(t23, o1, l19, j19);
and(u23, n1, l19, j19);
and(v23, m1, l19, j19);
and(w23, k1, m19, k19);
and(x23, y0, m19, t16);
and(y23, x0, m19, t16);
and(z23, w0, m19, t16);
and(a24, v0, m19, t16);
and(b24, u0, l19, s16);
and(c24, t0, l19, s16);
and(d24, s0, l19, s16);
and(e24, r0, l19, s16);
and(f24, p0, m19, t16);
and(g24, o0, w16, k19);
and(h24, n0, w16, k19);
and(i24, m0, w16, k19);
and(j24, l0, w16, k19);
and(k24, k0, v16, j19);
and(l24, j0, v16, j19);
and(m24, i0, v16, j19);
and(n24, h0, v16, j19);
and(o24, g0, v16, j19);
and(p24, e0, w16, k19);
and(q24, a0, k20);
and(r24, z, k20);
and(s24, y, l20);
and(t24, x, l20);
and(u24, v, k20);
and(v24, u, k20);
and(w24, t, l20);
and(x24, s, l20);
and(y24, r, m20);
and(z24, q, m20);
and(a25, p, m20);
and(b25, o, m20);
and(c25, n, n20);
and(d25, m, n20);
or(e25, f17, o20);
and(f25, f, m20);
and(g25, e, n20);
and(h25, d, n20);
not(t_68, l17);
not(t_69, u20);
or(i25, t_68, t_69);
not(t_70, m17);
not(t_71, v20);
or(j25, t_70, t_71);
not(k25, w20);
buf(l25, x20);
buf(m25, x20);
not(n25, y20);
not(o25, z20);
not(p25, a21);
or(q25, x17, b21, d21, c21);
not(t_72, e21);
not(t_73, f21);
or(r25, t_72, t_73);
not(t_74, h21);
not(t_75, j21);
or(s25, t_74, t_75);
not(t_76, l21);
not(t_77, n21);
or(t25, t_76, t_77);
not(t_78, q21);
not(t_79, s21);
or(u25, t_78, t_79);
not(t_80, u21);
not(t_81, w21);
or(v25, t_80, t_81);
not(t_82, y21);
not(t_83, a22);
or(w25, t_82, t_83);
not(t_84, c22);
not(t_85, e22);
or(x25, t_84, t_85);
not(t_86, h22);
not(t_87, j22);
or(y25, t_86, t_87);
not(z25, l22);
or(a26, n19, v22, e23, m22);
or(b26, o19, w22, f23, n22);
or(c26, p19, x22, g23, o22);
or(d26, q19, y22, h23, p22);
or(e26, r19, z22, i23, q22);
or(f26, s19, a23, j23, r22);
or(g26, t19, b23, k23, s22);
or(h26, u19, c23, l23, t22);
or(i26, v19, d23, m23, u22);
or(j26, w19, x23, g24, n23);
or(k26, x19, y23, h24, o23);
or(l26, y19, z23, i24, p23);
or(m26, z19, a24, j24, q23);
or(n26, a20, b24, k24, r23);
or(o26, b20, c24, l24, s23);
or(p26, c20, k22, m24, t23);
or(q26, d20, d24, n24, u23);
or(r26, e20, e24, o24, v23);
or(s26, f20, f24, p24, w23);
not(t26, i25);
not(u26, j25);
not(t_88, k25);
not(t_89, y25);
or(v26, t_88, t_89);
and(w26, n25, o25, l25);
not(x26, l25);
not(y26, m25);
and(z26, y20, z20, m25);
and(w11, p25, z25);
buf(b27, q25);
not(t_90, q25);
not(t_91, d15);
or(c27, t_90, t_91);
not(d27, r25);
not(t_92, h26);
not(t_93, f15);
or(e27, t_92, t_93);
buf(f27, s25);
buf(g27, s25);
not(h27, t25);
not(i27, u25);
not(j27, v25);
buf(k27, w25);
buf(l27, w25);
not(m27, x25);
and(n27, e26, k16);
not(o27, y25);
and(p27, s26, p16);
and(q27, k26, p16);
and(r27, n26, q6);
and(s27, s26, p6);
and(t27, k26, p6);
and(u27, j26, p6);
not(v27, a26);
buf(w27, b26);
buf(x27, c26);
buf(y27, c26);
buf(z27, d26);
buf(a28, e26);
not(b28, f26);
buf(c28, f26);
buf(d28, g26);
buf(e28, h26);
buf(f28, i26);
buf(g28, j26);
not(h28, j26);
not(i28, k26);
not(j28, k26);
buf(g12, l26);
buf(h12, m26);
buf(i12, n26);
buf(j12, o26);
buf(k12, p26);
buf(l12, q26);
buf(m12, r26);
not(r28, s26);
buf(s28, s26);
and(t28, g26, b17);
and(u28, f26, b17);
and(v28, e26, b17);
and(w28, h26, b17);
and(x28, i26, c17);
and(y28, d26, c17);
and(z28, c26, c17);
and(a29, b26, c17);
and(b29, p26, d17);
and(c29, o26, d17);
and(d29, n26, d17);
and(e29, r26, d17);
and(f29, q26, d17);
and(g29, s26, e17);
and(h29, m26, e17);
and(i29, l26, e17);
and(j29, k26, e17);
and(k29, t25, i25, g27);
and(l29, h27, t26, f27);
and(m29, x25, j25, l27);
and(n29, m27, u26, k27);
not(t_94, o27);
not(t_95, w20);
or(o29, t_94, t_95);
and(p29, o25, y20, y26);
and(q29, z20, n25, x26);
and(r29, c27, q25);
not(s29, b27);
and(t29, d15, c27);
and(u29, f15, e27);
not(v29, f27);
not(w29, g27);
not(t_96, j27);
not(t_97, u25);
or(x29, t_96, t_97);
not(t_98, i27);
not(t_99, v25);
or(y29, t_98, t_99);
not(z29, k27);
not(a30, l27);
not(b30, n27);
and(c30, g28, p16);
and(d30, g12, p16);
and(e30, h12, q6);
not(t_100, j28);
not(t_101, u16);
or(f30, t_100, t_101);
and(g30, r16, j6, w11, t20);
not(t_102, v27);
not(t_103, f28);
or(h30, t_102, t_103);
not(i30, w27);
not(j30, y27);
not(k30, z27);
not(l30, a28);
not(m30, c28);
not(n30, d28);
and(o30, e27, h26);
not(p30, e28);
not(q30, f28);
buf(r30, g28);
buf(s30, h28);
buf(t30, h28);
buf(u30, i28);
buf(v30, i28);
buf(w30, i28);
buf(x30, i28);
not(y30, j28);
not(z30, g12);
not(a31, h12);
not(b31, i12);
not(c31, j12);
not(d31, k12);
not(e31, l12);
not(f31, m12);
buf(g31, r28);
buf(h31, r28);
not(i31, s28);
and(j31, b28, n27, d0);
and(k31, r16, j6, b0, w11);
or(l31, t28, q24);
or(m31, u28, r24);
or(n31, y28, s24);
or(o31, a29, t24);
or(p31, w28, u24);
or(q31, v28, v24);
or(r31, z28, w24);
or(s31, x28, x24);
or(t31, e29, y24);
or(u31, b29, z24);
or(v31, c29, a25);
or(w31, d29, b25);
or(x31, i29, c25);
or(y31, g29, d25);
or(z31, f29, f25);
or(a32, h29, g25);
or(b32, j29, h25);
and(c32, i25, h27, v29);
and(d32, j25, m27, z29);
not(t_104, v26);
not(t_105, o29);
or(e32, t_104, t_105);
not(t_106, q29);
not(t_107, w26);
and(f32, t_106, t_107);
not(t_108, p29);
not(t_109, z26);
and(g32, t_108, t_109);
or(h32, r29, t29);
not(t_110, p30);
not(t_111, b27);
or(i32, t_110, t_111);
or(j32, o30, u29);
not(t_112, g21);
not(t_113, l31);
or(k32, t_112, t_113);
not(t_114, i21);
not(t_115, m31);
or(l32, t_114, t_115);
not(t_116, k21);
not(t_117, q31);
or(m32, t_116, t_117);
and(n32, t26, t25, w29);
not(t_118, m21);
not(t_119, n31);
or(o32, t_118, t_119);
not(t_120, o21);
not(t_121, r31);
or(p32, t_120, t_121);
not(t_122, p21);
not(t_123, o31);
or(q32, t_122, t_123);
not(t_124, x29);
not(t_125, y29);
or(r32, t_124, t_125);
not(t_126, r21);
not(t_127, s31);
or(s32, t_126, t_127);
not(t_128, t21);
not(t_129, t31);
or(t32, t_128, t_129);
not(t_130, v21);
not(t_131, z31);
or(u32, t_130, t_131);
not(t_132, x21);
not(t_133, u31);
or(v32, t_132, t_133);
not(t_134, z21);
not(t_135, v31);
or(w32, t_134, t_135);
not(t_136, b22);
not(t_137, w31);
or(x32, t_136, t_137);
and(y32, u26, x25, a30);
not(t_138, d22);
not(t_139, a32);
or(z32, t_138, t_139);
not(t_140, f22);
not(t_141, x31);
or(a33, t_140, t_141);
not(t_142, g22);
not(t_143, b32);
or(b33, t_142, t_143);
not(t_144, i22);
not(t_145, y31);
or(c33, t_144, t_145);
or(d33, e30, q27);
or(e33, r27, d30);
and(f33, f30, q6);
and(g33, f30, q16);
not(h33, f30);
buf(i33, f30);
not(t_146, q30);
not(t_147, a26);
or(j33, t_146, t_147);
not(t_148, j30);
not(t_149, w27);
or(k33, t_148, t_149);
not(t_150, i30);
not(t_151, y27);
or(l33, t_150, t_151);
not(t_152, l30);
not(t_153, z27);
or(m33, t_152, t_153);
not(t_154, k30);
not(t_155, a28);
or(n33, t_154, t_155);
not(t_156, n30);
not(t_157, c28);
or(o33, t_156, t_157);
not(t_158, m30);
not(t_159, d28);
or(p33, t_158, t_159);
not(t_160, s29);
not(t_161, e28);
or(q33, t_160, t_161);
not(r33, r30);
not(s33, s30);
not(t33, t30);
not(u33, u30);
not(v33, v30);
not(w33, w30);
not(x33, x30);
not(y33, y30);
not(t_162, i31);
not(t_163, y30);
or(z33, t_162, t_163);
buf(a34, z30);
buf(b34, z30);
buf(c34, z30);
buf(d34, z30);
buf(e34, a31);
buf(f34, a31);
buf(g34, a31);
not(h34, b31);
buf(i34, c31);
buf(j34, c31);
buf(k34, d31);
buf(l34, d31);
buf(m34, e31);
buf(n34, e31);
buf(o34, f31);
buf(p34, f31);
not(q34, g31);
not(r34, h31);
and(s34, d0, b28, b30);
buf(t34, j31);
not(u34, j31);
not(v34, j31);
buf(w34, j31);
not(x34, j31);
not(y34, l31);
not(z34, m31);
not(a35, n31);
not(b35, o31);
not(c35, q31);
not(d35, r31);
not(e35, s31);
not(f35, t31);
not(g35, u31);
not(h35, v31);
not(i35, w31);
not(j35, x31);
not(k35, y31);
not(l35, z31);
not(m35, a32);
not(n35, b32);
not(t_164, n32);
not(t_165, k29);
and(o35, t_164, t_165);
not(t_166, c32);
not(t_167, l29);
and(p35, t_166, t_167);
not(t_168, y32);
not(t_169, m29);
and(q35, t_168, t_169);
not(t_170, d32);
not(t_171, n29);
and(r35, t_170, t_171);
not(s35, e32);
not(t_172, g32);
not(t_173, f32);
or(t35, t_172, t_173);
not(u35, h32);
not(t_174, i32);
not(t_175, q33);
or(v35, t_174, t_175);
not(w35, j32);
not(t_176, y34);
not(t_177, d18);
or(x35, t_176, t_177);
not(t_178, z34);
not(t_179, f18);
or(y35, t_178, t_179);
not(t_180, c35);
not(t_181, h18);
or(z35, t_180, t_181);
not(t_182, a35);
not(t_183, j18);
or(a36, t_182, t_183);
not(t_184, d35);
not(t_185, l18);
or(b36, t_184, t_185);
not(t_186, b35);
not(t_187, n18);
or(c36, t_186, t_187);
not(d36, r32);
not(t_188, e35);
not(t_189, p18);
or(e36, t_188, t_189);
not(t_190, f35);
not(t_191, r18);
or(f36, t_190, t_191);
not(t_192, l35);
not(t_193, t18);
or(g36, t_192, t_193);
not(t_194, g35);
not(t_195, v18);
or(h36, t_194, t_195);
not(t_196, h35);
not(t_197, x18);
or(i36, t_196, t_197);
not(t_198, i35);
not(t_199, z18);
or(j36, t_198, t_199);
not(t_200, m35);
not(t_201, b19);
or(k36, t_200, t_201);
not(t_202, j35);
not(t_203, d19);
or(l36, t_202, t_203);
not(t_204, n35);
not(t_205, f19);
or(m36, t_204, t_205);
not(t_206, k35);
not(t_207, h19);
or(n36, t_206, t_207);
or(o36, f33, p27);
not(p36, h33);
not(q36, i33);
not(t_208, h30);
not(t_209, j33);
or(r36, t_208, t_209);
and(s36, b26, v34);
and(t36, b26, u34);
not(t_210, l33);
not(t_211, k33);
or(u36, t_210, t_211);
and(v36, x27, v34);
and(w36, x27, u34);
not(t_212, n33);
not(t_213, m33);
or(x36, t_212, t_213);
not(t_214, p33);
not(t_215, o33);
or(y36, t_214, t_215);
and(z36, i26, v34);
and(a37, i26, u34);
not(t_216, q34);
not(t_217, s30);
or(b37, t_216, t_217);
not(t_218, r34);
not(t_219, t30);
or(c37, t_218, t_219);
not(t_220, v33);
not(t_221, b34);
or(d37, t_220, t_221);
not(t_222, x33);
not(t_223, d34);
or(e37, t_222, t_223);
not(f37, a34);
not(g37, b34);
not(h37, c34);
not(i37, d34);
not(j37, e34);
not(k37, f34);
not(t_224, h34);
not(t_225, g34);
or(l37, t_224, t_225);
not(m37, g34);
and(n37, i12, w34);
and(o37, i12, t34);
and(p37, j12, w34);
and(q37, j12, t34);
not(r37, i34);
not(s37, j34);
not(t37, k34);
not(u37, l34);
not(v37, m34);
not(w37, n34);
and(x37, m12, v34);
and(y37, m12, u34);
not(z37, o34);
not(a38, p34);
not(t_226, s33);
not(t_227, g31);
or(b38, t_226, t_227);
not(t_228, t33);
not(t_229, h31);
or(c38, t_228, t_229);
not(t_230, y33);
not(t_231, s28);
or(d38, t_230, t_231);
buf(e38, s34);
buf(f38, s34);
not(g38, t34);
not(h38, w34);
buf(i38, x34);
buf(j38, x34);
not(t_232, o35);
not(t_233, p35);
or(k38, t_232, t_233);
not(t_234, q35);
not(t_235, r35);
or(l38, t_234, t_235);
not(t_236, s35);
not(t_237, t35);
or(m38, t_236, t_237);
not(n38, t35);
and(o38, h32, u35);
not(p38, v35);
and(q38, j32, w35);
not(t_238, x35);
not(t_239, k32);
or(r38, t_238, t_239);
not(t_240, y35);
not(t_241, l32);
or(s38, t_240, t_241);
not(t_242, z35);
not(t_243, m32);
or(t38, t_242, t_243);
not(t_244, a36);
not(t_245, o32);
or(u38, t_244, t_245);
not(t_246, b36);
not(t_247, p32);
or(v38, t_246, t_247);
not(t_248, c36);
not(t_249, q32);
or(w38, t_248, t_249);
not(t_250, e36);
not(t_251, s32);
or(x38, t_250, t_251);
not(t_252, f36);
not(t_253, t32);
or(y38, t_252, t_253);
not(t_254, g36);
not(t_255, u32);
or(z38, t_254, t_255);
not(t_256, h36);
not(t_257, v32);
or(a39, t_256, t_257);
not(t_258, i36);
not(t_259, w32);
or(b39, t_258, t_259);
not(t_260, j36);
not(t_261, x32);
or(c39, t_260, t_261);
not(t_262, k36);
not(t_263, z32);
or(d39, t_262, t_263);
not(t_264, l36);
not(t_265, a33);
or(e39, t_264, t_265);
not(t_266, m36);
not(t_267, b33);
or(f39, t_266, t_267);
not(t_268, n36);
not(t_269, c33);
or(g39, t_268, t_269);
not(h39, r36);
not(i39, u36);
buf(j39, x36);
buf(k39, x36);
not(l39, y36);
not(t_270, b38);
not(t_271, b37);
or(m39, t_270, t_271);
not(t_272, c38);
not(t_273, c37);
or(n39, t_272, t_273);
not(t_274, g37);
not(t_275, v30);
or(o39, t_274, t_275);
not(t_276, i37);
not(t_277, x30);
or(p39, t_276, t_277);
not(t_278, z33);
not(t_279, d38);
or(q39, t_278, t_279);
and(r39, i12, h38);
and(s39, i12, g38);
not(t_280, m37);
not(t_281, b31);
or(t39, t_280, t_281);
and(u39, j12, h38);
and(v39, j12, g38);
not(t_282, t37);
not(t_283, i34);
or(w39, t_282, t_283);
not(t_284, u37);
not(t_285, j34);
or(x39, t_284, t_285);
and(y39, k12, h38);
and(z39, k12, g38);
not(t_286, r37);
not(t_287, k34);
or(a40, t_286, t_287);
not(t_288, s37);
not(t_289, l34);
or(b40, t_288, t_289);
and(c40, l12, h38);
and(d40, l12, g38);
not(t_290, z37);
not(t_291, m34);
or(e40, t_290, t_291);
not(t_292, a38);
not(t_293, n34);
or(f40, t_292, t_293);
not(t_294, v37);
not(t_295, o34);
or(g40, t_294, t_295);
not(t_296, w37);
not(t_297, p34);
or(h40, t_296, t_297);
buf(i40, e38);
buf(j40, e38);
buf(k40, f38);
buf(l40, f38);
buf(m40, i38);
buf(n40, i38);
buf(o40, i38);
buf(p40, j38);
buf(q40, j38);
buf(r40, j38);
not(s40, k38);
not(t40, l38);
not(t_298, n38);
not(t_299, e32);
or(u40, t_298, t_299);
or(v40, u35, o38);
not(t_300, l39);
not(t_301, v35);
or(w40, t_300, t_301);
not(t_302, d27);
not(t_303, k38);
or(x40, t_302, t_303);
or(y40, w35, q38);
not(z40, r38);
not(a41, s38);
not(b41, t38);
not(c41, u38);
and(d41, q15, n40);
and(e41, q15, q40);
not(f41, v38);
and(g41, s15, n40);
and(h41, s15, q40);
not(i41, w38);
not(t_304, d36);
not(t_305, l38);
or(j41, t_304, t_305);
and(k41, u15, n40);
and(l41, u15, q40);
not(m41, x38);
and(n41, w15, n40);
and(o41, w15, q40);
not(p41, y38);
and(q41, y15, m40);
and(r41, y15, p40);
not(s41, z38);
and(t41, a16, m40);
and(u41, a16, p40);
not(v41, a39);
and(w41, c16, m40);
and(x41, c16, p40);
not(y41, b39);
and(z41, e16, m40);
and(a42, e16, p40);
not(b42, c39);
and(c42, g16, o40);
and(d42, g16, r40);
not(e42, d39);
and(f42, i16, o40);
and(g42, i16, r40);
not(h42, e39);
and(i42, l16, r40);
and(j42, l16, o40);
not(k42, f39);
and(l42, n16, o40);
and(m42, n16, r40);
not(n42, g39);
not(t_306, p36);
not(t_307, q39);
or(o42, t_306, t_307);
and(p42, u36, r36, k39);
and(q42, i39, h39, j39);
and(r42, s36, i40);
and(s42, t36, j40);
and(t42, v36, i40);
and(u42, w36, j40);
not(v42, j39);
not(w42, k39);
not(t_308, p38);
not(t_309, y36);
or(x42, t_308, t_309);
and(y42, z36, i40);
and(z42, a37, j40);
not(a43, m39);
not(b43, n39);
not(t_310, d37);
not(t_311, o39);
or(c43, t_310, t_311);
not(t_312, e37);
not(t_313, p39);
or(d43, t_312, t_313);
not(e43, q39);
not(t_314, t39);
not(t_315, l37);
or(f43, t_314, t_315);
or(g43, n37, r39);
or(h43, o37, s39);
or(i43, p37, u39);
or(j43, q37, v39);
not(t_316, a40);
not(t_317, w39);
or(k43, t_316, t_317);
not(t_318, b40);
not(t_319, x39);
or(l43, t_318, t_319);
not(t_320, g40);
not(t_321, e40);
or(m43, t_320, t_321);
not(t_322, h40);
not(t_323, f40);
or(n43, t_322, t_323);
and(o43, x37, i40);
and(p43, y37, j40);
not(q43, m40);
not(r43, o40);
not(s43, p40);
not(t43, r40);
and(u43, y39, r20);
and(v43, c40, r20);
and(w43, z39, s20);
and(x43, d40, s20);
not(t_324, m38);
not(t_325, u40);
or(y43, t_324, t_325);
not(t_326, w40);
not(t_327, x42);
or(z43, t_326, t_327);
not(t_328, s40);
not(t_329, r25);
or(a44, t_328, t_329);
and(b44, h15, q43);
and(c44, h15, s43);
and(d44, j15, q43);
and(e44, j15, s43);
and(f44, a41, b41, c41, f41, i41);
and(g44, l15, r43);
and(h44, l15, t43);
and(i44, n15, r43);
and(j44, n15, t43);
and(k44, q15, r43);
and(l44, q15, t43);
and(m44, s15, r43);
and(n44, s15, t43);
not(t_330, t40);
not(t_331, r32);
or(o44, t_330, t_331);
and(p44, m41, p41, s41, v41, y41);
and(q44, b42, e42, h42, k42, n42);
not(t_332, e43);
not(t_333, h33);
or(r44, t_332, t_333);
and(s44, r36, i39, v42);
not(t44, r42);
not(u44, s42);
and(v44, h39, u36, w42);
not(w44, t42);
not(x44, u42);
not(y44, y42);
not(z44, z42);
not(a45, c43);
buf(b45, d43);
buf(c45, d43);
buf(d45, f43);
buf(e45, f43);
not(f45, k43);
not(g45, l43);
not(h45, m43);
not(i45, n43);
not(j45, o43);
not(k45, p43);
and(l45, g41, k40);
and(m45, k41, k40);
and(n45, n41, k40);
and(o45, d41, k40);
and(p45, h41, l40);
and(q45, l41, l40);
and(r45, o41, l40);
and(s45, e41, l40);
and(t45, p31, z40);
and(u45, q41, p20);
and(v45, t41, p20);
and(w45, r41, q20);
and(x45, u41, q20);
and(y45, g43, r20);
and(z45, i43, r20);
not(a46, u43);
not(b46, v43);
and(c46, h43, s20);
and(d46, j43, s20);
not(e46, w43);
not(f46, x43);
not(g46, y43);
not(h46, z43);
not(t_334, x40);
not(t_335, a44);
or(i46, t_334, t_335);
and(j46, t45, f44);
not(t_336, j41);
not(t_337, o44);
or(k46, t_336, t_337);
and(l46, p44, q44);
or(m46, w41, b44);
or(n46, x41, c44);
or(o46, z41, d44);
or(p46, a42, e44);
or(q46, c42, g44);
or(r46, d42, h44);
or(s46, f42, i44);
or(t46, g42, j44);
or(u46, i42, l44);
or(v46, j42, k44);
or(w46, l42, m44);
or(x46, m42, n44);
not(t_338, r44);
not(t_339, o42);
or(y46, t_338, t_339);
and(z46, n39, i33, b45);
and(a47, b43, q36, c45);
not(t_340, v44);
not(t_341, p42);
and(b47, t_340, t_341);
not(t_342, s44);
not(t_343, q42);
and(c47, t_342, t_343);
and(d47, l45, t44);
buf(e47, t44);
and(f47, p45, u44);
buf(g47, u44);
and(h47, o45, w44);
buf(i47, w44);
and(j47, s45, x44);
buf(k47, x44);
and(l47, m45, y44);
buf(m47, y44);
and(n47, q45, z44);
buf(o47, z44);
and(p47, c43, m39, e45);
and(q47, a45, a43, d45);
not(r47, b45);
not(s47, c45);
not(t47, d45);
not(u47, e45);
not(t_344, h45);
not(t_345, k43);
or(v47, t_344, t_345);
not(t_346, i45);
not(t_347, l43);
or(w47, t_346, t_347);
not(t_348, f45);
not(t_349, m43);
or(x47, t_348, t_349);
not(t_350, g45);
not(t_351, n43);
or(y47, t_350, t_351);
and(z47, j45, n45);
buf(a48, j45);
and(b48, k45, r45);
buf(c48, k45);
buf(d48, l45);
buf(e48, m45);
buf(f48, n45);
buf(g48, o45);
buf(h48, p45);
buf(i48, q45);
buf(j48, r45);
buf(k48, s45);
and(l48, u45, b46);
buf(m48, u45);
and(n48, v45, a46);
buf(o48, v45);
and(p48, w45, f46);
buf(q48, w45);
and(r48, x45, e46);
buf(s48, x45);
not(t48, y45);
not(u48, z45);
buf(v48, a46);
buf(w48, b46);
not(x48, c46);
not(y48, d46);
buf(z48, e46);
buf(a49, f46);
buf(b49, q46);
buf(c49, r46);
buf(d49, s46);
buf(e49, t46);
buf(f49, u46);
buf(g49, v46);
not(h49, y46);
and(i49, i33, b43, s47);
and(j49, q36, n39, r47);
not(t_352, b47);
not(t_353, c47);
or(k49, t_352, t_353);
not(l49, e47);
not(m49, g47);
not(n49, i47);
not(o49, k47);
not(p49, m47);
not(q49, o47);
not(t_354, r33);
not(t_355, y46);
or(r49, t_354, t_355);
and(s49, m39, a45, t47);
and(t49, a43, c43, u47);
and(u49, v46, i28);
and(v49, u46, i28);
and(w49, s46, z30);
and(x49, t46, z30);
and(y49, q46, a31);
and(z49, r46, a31);
not(t_356, x47);
not(t_357, v47);
or(a50, t_356, t_357);
not(t_358, y47);
not(t_359, w47);
or(b50, t_358, t_359);
not(c50, a48);
not(d50, c48);
and(e50, w46, r28);
and(f50, x46, r28);
not(g50, d48);
not(h50, e48);
not(i50, f48);
not(j50, g48);
not(k50, h48);
not(l50, i48);
not(m50, j48);
not(n50, k48);
and(v12, g46, j);
and(y12, l46, j46, e25);
not(q50, m48);
not(r50, o48);
and(s50, m46, p20);
and(t50, o46, p20);
not(u50, q48);
not(v50, s48);
and(w50, n46, q20);
and(x50, p46, q20);
buf(y50, t48);
buf(z50, u48);
not(a51, v48);
not(b51, w48);
buf(c51, x48);
buf(d51, y48);
not(e51, z48);
not(f51, a49);
not(t_360, h46);
not(t_361, k49);
or(g51, t_360, t_361);
not(h51, b49);
not(i51, c49);
not(j51, d49);
not(k51, e49);
not(l51, f49);
not(m51, g49);
not(t_362, j49);
not(t_363, z46);
and(n51, t_362, t_363);
not(t_364, i49);
not(t_365, a47);
and(o51, t_364, t_365);
not(p51, k49);
not(t_366, g50);
not(t_367, e47);
or(q51, t_366, t_367);
not(t_368, k50);
not(t_369, g47);
or(r51, t_368, t_369);
not(t_370, j50);
not(t_371, i47);
or(s51, t_370, t_371);
not(t_372, n50);
not(t_373, k47);
or(t51, t_372, t_373);
not(t_374, h50);
not(t_375, m47);
or(u51, t_374, t_375);
not(t_376, l50);
not(t_377, o47);
or(v51, t_376, t_377);
not(t_378, h49);
not(t_379, r30);
or(w51, t_378, t_379);
not(t_380, t49);
not(t_381, p47);
and(x51, t_380, t_381);
not(t_382, s49);
not(t_383, q47);
and(y51, t_382, t_383);
not(t_384, u33);
not(t_385, f49);
or(z51, t_384, t_385);
not(t_386, w33);
not(t_387, g49);
or(a52, t_386, t_387);
not(t_388, f37);
not(t_389, e49);
or(b52, t_388, t_389);
not(t_390, h37);
not(t_391, d49);
or(c52, t_390, t_391);
not(t_392, j37);
not(t_393, c49);
or(d52, t_392, t_393);
not(t_394, k37);
not(t_395, b49);
or(e52, t_394, t_395);
not(f52, a50);
not(g52, b50);
not(t_396, i50);
not(t_397, a48);
or(h52, t_396, t_397);
not(t_398, m50);
not(t_399, c48);
or(i52, t_398, t_399);
not(t_400, l49);
not(t_401, d48);
or(j52, t_400, t_401);
not(t_402, p49);
not(t_403, e48);
or(k52, t_402, t_403);
not(t_404, c50);
not(t_405, f48);
or(l52, t_404, t_405);
not(t_406, n49);
not(t_407, g48);
or(m52, t_406, t_407);
not(t_408, m49);
not(t_409, h48);
or(n52, t_408, t_409);
not(t_410, q49);
not(t_411, i48);
or(o52, t_410, t_411);
not(t_412, d50);
not(t_413, j48);
or(p52, t_412, t_413);
not(t_414, o49);
not(t_415, k48);
or(q52, t_414, t_415);
not(r52, v12);
not(t_416, b51);
not(t_417, m48);
or(s52, t_416, t_417);
not(t_418, a51);
not(t_419, o48);
or(t52, t_418, t_419);
buf(u52, s50);
buf(v52, t50);
not(t_420, f51);
not(t_421, q48);
or(w52, t_420, t_421);
not(t_422, e51);
not(t_423, s48);
or(x52, t_422, t_423);
buf(y52, w50);
buf(z52, x50);
not(a53, y50);
and(b53, t50, t48);
and(c53, s50, u48);
not(d53, z50);
not(t_424, r50);
not(t_425, v48);
or(e53, t_424, t_425);
not(t_426, q50);
not(t_427, w48);
or(f53, t_426, t_427);
not(g53, c51);
and(h53, x50, x48);
and(i53, w50, y48);
not(j53, d51);
not(t_428, v50);
not(t_429, z48);
or(k53, t_428, t_429);
not(t_430, u50);
not(t_431, a49);
or(l53, t_430, t_431);
not(t_432, p51);
not(t_433, z43);
or(m53, t_432, t_433);
not(t_434, n51);
not(t_435, o51);
or(n53, t_434, t_435);
not(t_436, j52);
not(t_437, q51);
or(o53, t_436, t_437);
not(t_438, n52);
not(t_439, r51);
or(p53, t_438, t_439);
not(t_440, m52);
not(t_441, s51);
or(q53, t_440, t_441);
not(t_442, q52);
not(t_443, t51);
or(r53, t_442, t_443);
not(t_444, k52);
not(t_445, u51);
or(s53, t_444, t_445);
not(t_446, o52);
not(t_447, v51);
or(t53, t_446, t_447);
not(t_448, w51);
not(t_449, r49);
or(u53, t_448, t_449);
not(t_450, x51);
not(t_451, y51);
or(v53, t_450, t_451);
not(t_452, l51);
not(t_453, u30);
or(w53, t_452, t_453);
not(t_454, m51);
not(t_455, w30);
or(x53, t_454, t_455);
not(t_456, k51);
not(t_457, a34);
or(y53, t_456, t_457);
not(t_458, j51);
not(t_459, c34);
or(z53, t_458, t_459);
not(t_460, i51);
not(t_461, e34);
or(a54, t_460, t_461);
not(t_462, h51);
not(t_463, f34);
or(b54, t_462, t_463);
not(t_464, l52);
not(t_465, h52);
or(c54, t_464, t_465);
not(t_466, p52);
not(t_467, i52);
or(d54, t_466, t_467);
not(t_468, s52);
not(t_469, f53);
or(e54, t_468, t_469);
not(t_470, t52);
not(t_471, e53);
or(f54, t_470, t_471);
not(t_472, d53);
not(t_473, u52);
or(g54, t_472, t_473);
not(h54, u52);
not(t_474, a53);
not(t_475, v52);
or(i54, t_474, t_475);
not(j54, v52);
not(t_476, w52);
not(t_477, l53);
or(k54, t_476, t_477);
not(t_478, x52);
not(t_479, k53);
or(l54, t_478, t_479);
not(t_480, j53);
not(t_481, y52);
or(m54, t_480, t_481);
not(n54, y52);
not(t_482, g53);
not(t_483, z52);
or(o54, t_482, t_483);
not(p54, z52);
not(t_484, g51);
not(t_485, m53);
or(q54, t_484, t_485);
and(r54, u53, q16);
not(s54, n53);
and(t54, q53, d47);
and(u54, o53, c54, s53, q53);
and(v54, r53, f47);
and(w54, p53, d54, t53, r53);
and(x54, o53, q53, l47);
and(y54, p53, r53, n47);
not(z54, v53);
not(t_486, z51);
not(t_487, w53);
or(a55, t_486, t_487);
not(t_488, a52);
not(t_489, x53);
or(b55, t_488, t_489);
not(t_490, b52);
not(t_491, y53);
or(c55, t_490, t_491);
not(t_492, c52);
not(t_493, z53);
or(d55, t_492, t_493);
not(t_494, d52);
not(t_495, a54);
or(e55, t_494, t_495);
not(t_496, e52);
not(t_497, b54);
or(f55, t_496, t_497);
not(t_498, f52);
not(t_499, v53);
or(g55, t_498, t_499);
not(t_500, g52);
not(t_501, n53);
or(h55, t_500, t_501);
and(i55, s53, q53, z47, o53);
and(j55, t53, r53, b48, p53);
and(k55, e54, n48);
and(l55, k54, r48);
not(t_502, j54);
not(t_503, y50);
or(m55, t_502, t_503);
and(n55, f54, e54, c53);
not(t_504, h54);
not(t_505, z50);
or(o55, t_504, t_505);
not(t_506, p54);
not(t_507, c51);
or(p55, t_506, t_507);
and(q55, l54, k54, i53);
not(t_508, n54);
not(t_509, d51);
or(r55, t_508, t_509);
not(s55, q54);
not(t55, u54);
not(u55, w54);
or(v55, i55, x54, t54, h47);
or(w55, j55, y54, v54, j47);
and(x55, d55, u49);
and(y55, c55, v49);
not(t_510, z54);
not(t_511, a50);
or(z55, t_510, t_511);
not(t_512, s54);
not(t_513, b50);
or(a56, t_512, t_513);
and(b56, b55, d55, e50);
and(c56, a55, c55, f50);
not(t_514, g54);
not(t_515, o55);
or(d56, t_514, t_515);
not(t_516, i54);
not(t_517, m55);
or(e56, t_516, t_517);
not(t_518, m54);
not(t_519, r55);
or(f56, t_518, t_519);
not(t_520, o54);
not(t_521, p55);
or(g56, t_520, t_521);
not(h56, v55);
not(i56, w55);
or(j56, b56, x55, w49);
or(k56, c56, y55, x49);
and(l56, e56, d56, e54, y49, f54);
and(m56, g56, f56, k54, z49, l54);
not(t_522, g55);
not(t_523, z55);
or(n56, t_522, t_523);
not(t_524, h55);
not(t_525, a56);
or(o56, t_524, t_525);
and(b13, s55, j20);
and(q56, f54, f55, d56, e54, e56);
and(r56, l54, e55, f56, k54, g56);
and(s56, d56, e54, b53, f54);
and(t56, f56, k54, h53, l54);
and(u56, o56, q6);
not(t_526, t55);
not(t_527, h56);
or(v56, t_526, t_527);
not(t_528, u55);
not(t_529, i56);
or(w56, t_528, t_529);
and(x56, q56, j56);
and(y56, r56, k56);
not(z56, n56);
not(a57, b13);
or(b57, l56, s56, n55, k55, l48);
or(c57, m56, t56, q55, l55, p48);
or(d57, u56, c30);
or(e57, x56, b57);
or(f57, y56, c57);
and(e13, z56, j20);
and(h57, v56, e57);
and(i57, w56, f57);
not(j57, e57);
not(k57, f57);
not(l57, e13);
and(m57, a57, l57, i46);
and(n57, v55, j57);
and(o57, w55, k57);
or(p57, h57, n57);
or(f13, i57, o57);
not(t_530, p57);
not(t_531, f13);
or(r57, t_530, t_531);
and(s57, r57, p57);
and(t57, f13, r57);
or(u57, s57, t57);
not(v57, u57);
and(w57, u57, v57);
or(x57, v57, w57);
and(y57, k46, r52, x57);
and(h13, m57, y57, w11);
buf(z7, k3);
buf(a8, l3);
buf(b8, m3);
buf(c8, n3);
buf(d8, o3);
buf(e8, p3);
buf(f8, q3);
buf(g8, r3);
buf(h8, s3);
buf(i8, t3);
buf(j8, u3);
buf(k8, v3);
buf(l8, w3);
buf(m8, x3);
buf(n8, y3);
buf(o8, z3);
buf(p8, a4);
buf(q8, b4);
buf(r8, c4);
buf(s8, d4);
buf(t8, e4);
buf(u8, f4);
buf(v8, g4);
buf(w8, h4);
buf(x8, i4);
buf(y8, j4);
buf(z8, k4);
buf(a9, l4);
buf(b9, m4);
buf(c9, n4);
buf(d9, o4);
buf(e9, p4);
buf(f9, q4);
buf(g9, r4);
buf(h9, s4);
buf(i9, t4);
buf(j9, u4);
buf(k9, v4);
buf(l9, w4);
buf(m9, x4);
buf(n9, y4);
buf(o9, z4);
buf(p9, a5);
buf(q9, b5);
buf(r9, c5);
buf(s9, d5);
buf(t9, e5);
buf(u9, f5);
buf(v9, g5);
buf(w9, h5);
buf(x9, i5);
buf(y9, j5);
buf(z9, k5);
buf(a10, l5);
buf(b10, m5);
buf(c10, n5);
buf(d10, o5);
buf(e10, p5);
buf(f10, q5);
buf(g10, r5);
buf(h10, s5);
buf(i10, t5);
buf(j10, u5);
buf(k10, v5);
buf(l10, w5);
buf(m10, x5);
buf(n10, y5);
buf(o10, z5);
buf(p10, a6);
buf(q10, b6);
buf(r10, c6);
buf(s10, d6);
buf(t10, e6);
buf(u10, f6);
buf(v10, g6);
buf(w10, h6);
buf(x10, i6);
buf(y10, i6);
buf(z10, i6);
buf(a11, r6);
buf(b11, r6);
buf(c11, e7);
buf(d11, e7);
buf(e11, e7);
buf(n12, d33);
buf(o12, d33);
buf(p12, e33);
buf(q12, e33);
buf(s12, o36);
buf(t12, o36);
buf(c13, d57);
buf(d13, d57);
endmodule
module top;
	parameter in_width = 233,
		patterns = 5000,
		step = 1;
	reg [1:in_width] in_mem[1:patterns];
	integer index;

	wire i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,
		i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,
		i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,
		i30,i31,i32,i33,i34,i35,i36,i37,i38,i39,
		i40,i41,i42,i43,i44,i45,i46,i47,i48,i49,
		i50,i51,i52,i53,i54,i55,i56,i57,i58,i59,
		i60,i61,i62,i63,i64,i65,i66,i67,i68,i69,
		i70,i71,i72,i73,i74,i75,i76,i77,i78,i79,
		i80,i81,i82,i83,i84,i85,i86,i87,i88,i89,
		i90,i91,i92,i93,i94,i95,i96,i97,i98,i99,
		i100,i101,i102,i103,i104,i105,i106,i107,i108,i109,
		i110,i111,i112,i113,i114,i115,i116,i117,i118,i119,
		i120,i121,i122,i123,i124,i125,i126,i127,i128,i129,
		i130,i131,i132,i133,i134,i135,i136,i137,i138,i139,
		i140,i141,i142,i143,i144,i145,i146,i147,i148,i149,
		i150,i151,i152,i153,i154,i155,i156,i157,i158,i159,
		i160,i161,i162,i163,i164,i165,i166,i167,i168,i169,
		i170,i171,i172,i173,i174,i175,i176,i177,i178,i179,
		i180,i181,i182,i183,i184,i185,i186,i187,i188,i189,
		i190,i191,i192,i193,i194,i195,i196,i197,i198,i199,
		i200,i201,i202,i203,i204,i205,i206,i207,i208,i209,
		i210,i211,i212,i213,i214,i215,i216,i217,i218,i219,
		i220,i221,i222,i223,i224,i225,i226,i227,i228,i229,
		i230,i231,i232;

	assign {i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,
		i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,
		i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,
		i30,i31,i32,i33,i34,i35,i36,i37,i38,i39,
		i40,i41,i42,i43,i44,i45,i46,i47,i48,i49,
		i50,i51,i52,i53,i54,i55,i56,i57,i58,i59,
		i60,i61,i62,i63,i64,i65,i66,i67,i68,i69,
		i70,i71,i72,i73,i74,i75,i76,i77,i78,i79,
		i80,i81,i82,i83,i84,i85,i86,i87,i88,i89,
		i90,i91,i92,i93,i94,i95,i96,i97,i98,i99,
		i100,i101,i102,i103,i104,i105,i106,i107,i108,i109,
		i110,i111,i112,i113,i114,i115,i116,i117,i118,i119,
		i120,i121,i122,i123,i124,i125,i126,i127,i128,i129,
		i130,i131,i132,i133,i134,i135,i136,i137,i138,i139,
		i140,i141,i142,i143,i144,i145,i146,i147,i148,i149,
		i150,i151,i152,i153,i154,i155,i156,i157,i158,i159,
		i160,i161,i162,i163,i164,i165,i166,i167,i168,i169,
		i170,i171,i172,i173,i174,i175,i176,i177,i178,i179,
		i180,i181,i182,i183,i184,i185,i186,i187,i188,i189,
		i190,i191,i192,i193,i194,i195,i196,i197,i198,i199,
		i200,i201,i202,i203,i204,i205,i206,i207,i208,i209,
		i210,i211,i212,i213,i214,i215,i216,i217,i218,i219,
		i220,i221,i222,i223,i224,i225,i226,i227,i228,i229,
		i230,i231,i232} = 
		$getpattern(in_mem[index]);

	initial $monitor($time,,o0,o1,o2,o3,o4,o5,o6,o7,o8,o9,
		o10,o11,o12,o13,o14,o15,o16,o17,o18,o19,
		o20,o21,o22,o23,o24,o25,o26,o27,o28,o29,
		o30,o31,o32,o33,o34,o35,o36,o37,o38,o39,
		o40,o41,o42,o43,o44,o45,o46,o47,o48,o49,
		o50,o51,o52,o53,o54,o55,o56,o57,o58,o59,
		o60,o61,o62,o63,o64,o65,o66,o67,o68,o69,
		o70,o71,o72,o73,o74,o75,o76,o77,o78,o79,
		o80,o81,o82,o83,o84,o85,o86,o87,o88,o89,
		o90,o91,o92,o93,o94,o95,o96,o97,o98,o99,
		o100,o101,o102,o103,o104,o105,o106,o107,o108,o109,
		o110,o111,o112,o113,o114,o115,o116,o117,o118,o119,
		o120,o121,o122,o123,o124,o125,o126,o127,o128,o129,
		o130,o131,o132,o133,o134,o135,o136,o137,o138,o139);
	initial
		begin
			$readmemb("patt.mem", in_mem);
			for(index = 1; index <= patterns; index = index + 1)
				#step;
		end

	foobar cct(o0,o1,o2,o3,o4,o5,o6,o7,o8,o9,
		o10,o11,o12,o13,o14,o15,o16,o17,o18,o19,
		o20,o21,o22,o23,o24,o25,o26,o27,o28,o29,
		o30,o31,o32,o33,o34,o35,o36,o37,o38,o39,
		o40,o41,o42,o43,o44,o45,o46,o47,o48,o49,
		o50,o51,o52,o53,o54,o55,o56,o57,o58,o59,
		o60,o61,o62,o63,o64,o65,o66,o67,o68,o69,
		o70,o71,o72,o73,o74,o75,o76,o77,o78,o79,
		o80,o81,o82,o83,o84,o85,o86,o87,o88,o89,
		o90,o91,o92,o93,o94,o95,o96,o97,o98,o99,
		o100,o101,o102,o103,o104,o105,o106,o107,o108,o109,
		o110,o111,o112,o113,o114,o115,o116,o117,o118,o119,
		o120,o121,o122,o123,o124,o125,o126,o127,o128,o129,
		o130,o131,o132,o133,o134,o135,o136,o137,o138,o139,
		i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,
		i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,
		i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,
		i30,i31,i32,i33,i34,i35,i36,i37,i38,i39,
		i40,i41,i42,i43,i44,i45,i46,i47,i48,i49,
		i50,i51,i52,i53,i54,i55,i56,i57,i58,i59,
		i60,i61,i62,i63,i64,i65,i66,i67,i68,i69,
		i70,i71,i72,i73,i74,i75,i76,i77,i78,i79,
		i80,i81,i82,i83,i84,i85,i86,i87,i88,i89,
		i90,i91,i92,i93,i94,i95,i96,i97,i98,i99,
		i100,i101,i102,i103,i104,i105,i106,i107,i108,i109,
		i110,i111,i112,i113,i114,i115,i116,i117,i118,i119,
		i120,i121,i122,i123,i124,i125,i126,i127,i128,i129,
		i130,i131,i132,i133,i134,i135,i136,i137,i138,i139,
		i140,i141,i142,i143,i144,i145,i146,i147,i148,i149,
		i150,i151,i152,i153,i154,i155,i156,i157,i158,i159,
		i160,i161,i162,i163,i164,i165,i166,i167,i168,i169,
		i170,i171,i172,i173,i174,i175,i176,i177,i178,i179,
		i180,i181,i182,i183,i184,i185,i186,i187,i188,i189,
		i190,i191,i192,i193,i194,i195,i196,i197,i198,i199,
		i200,i201,i202,i203,i204,i205,i206,i207,i208,i209,
		i210,i211,i212,i213,i214,i215,i216,i217,i218,i219,
		i220,i221,i222,i223,i224,i225,i226,i227,i228,i229,
		i230,i231,i232);
endmodule