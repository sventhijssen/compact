// IWLS benchmark module "DES" printed on Wed May 29 16:08:42 2002
module DES(\data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , \reset<0> , \encrypt<0> , \load_key<0> , \inreg<55> , \inreg<54> , \inreg<53> , \inreg<52> , \inreg<51> , \inreg<50> , \inreg<49> , \inreg<48> , \inreg<47> , \inreg<46> , \inreg<45> , \inreg<44> , \inreg<43> , \inreg<42> , \inreg<41> , \inreg<40> , \inreg<39> , \inreg<38> , \inreg<37> , \inreg<36> , \inreg<35> , \inreg<34> , \inreg<33> , \inreg<32> , \inreg<31> , \inreg<30> , \inreg<29> , \inreg<28> , \inreg<27> , \inreg<26> , \inreg<25> , \inreg<24> , \inreg<23> , \inreg<22> , \inreg<21> , \inreg<20> , \inreg<19> , \inreg<18> , \inreg<17> , \inreg<16> , \inreg<15> , \inreg<14> , \inreg<13> , \inreg<12> , \inreg<11> , \inreg<10> , \inreg<9> , \inreg<8> , \inreg<7> , \inreg<6> , \inreg<5> , \inreg<4> , \inreg<3> , \inreg<2> , \inreg<1> , \inreg<0> , \outreg<63> , \outreg<62> , \outreg<61> , \outreg<60> , \outreg<59> , \outreg<58> , \outreg<57> , \outreg<56> , \outreg<55> , \outreg<54> , \outreg<53> , \outreg<52> , \outreg<51> , \outreg<50> , \outreg<49> , \outreg<48> , \outreg<47> , \outreg<46> , \outreg<45> , \outreg<44> , \outreg<43> , \outreg<42> , \outreg<41> , \outreg<40> , \outreg<39> , \outreg<38> , \outreg<37> , \outreg<36> , \outreg<35> , \outreg<34> , \outreg<33> , \outreg<32> , \outreg<31> , \outreg<30> , \outreg<29> , \outreg<28> , \outreg<27> , \outreg<26> , \outreg<25> , \outreg<24> , \outreg<23> , \outreg<22> , \outreg<21> , \outreg<20> , \outreg<19> , \outreg<18> , \outreg<17> , \outreg<16> , \outreg<15> , \outreg<14> , \outreg<13> , \outreg<12> , \outreg<11> , \outreg<10> , \outreg<9> , \outreg<8> , \outreg<7> , \outreg<6> , \outreg<5> , \outreg<4> , \outreg<3> , \outreg<2> , \outreg<1> , \outreg<0> , \data<63> , \data<62> , \data<61> , \data<60> , \data<59> , \data<58> , \data<57> , \data<56> , \data<55> , \data<54> , \data<53> , \data<52> , \data<51> , \data<50> , \data<49> , \data<48> , \data<47> , \data<46> , \data<45> , \data<44> , \data<43> , \data<42> , \data<41> , \data<40> , \data<39> , \data<38> , \data<37> , \data<36> , \data<35> , \data<34> , \data<33> , \data<32> , \data<31> , \data<30> , \data<29> , \data<28> , \data<27> , \data<26> , \data<25> , \data<24> , \data<23> , \data<22> , \data<21> , \data<20> , \data<19> , \data<18> , \data<17> , \data<16> , \data<15> , \data<14> , \data<13> , \data<12> , \data<11> , \data<10> , \data<9> , \data<8> , \data<7> , \data<6> , \data<5> , \data<4> , \data<3> , \data<2> , \data<1> , \data<0> , \count<3> , \count<2> , \count<1> , \count<0> , \C<27> , \C<26> , \C<25> , \C<24> , \C<23> , \C<22> , \C<21> , \C<20> , \C<19> , \C<18> , \C<17> , \C<16> , \C<15> , \C<14> , \C<13> , \C<12> , \C<11> , \C<10> , \C<9> , \C<8> , \C<7> , \C<6> , \C<5> , \C<4> , \C<3> , \C<2> , \C<1> , \C<0> , \D<27> , \D<26> , \D<25> , \D<24> , \D<23> , \D<22> , \D<21> , \D<20> , \D<19> , \D<18> , \D<17> , \D<16> , \D<15> , \D<14> , \D<13> , \D<12> , \D<11> , \D<10> , \D<9> , \D<8> , \D<7> , \D<6> , \D<5> , \D<4> , \D<3> , \D<2> , \D<1> , \D<0> , \encrypt_mode<0> , \inreg_new<55> , \inreg_new<54> , \inreg_new<53> , \inreg_new<52> , \inreg_new<51> , \inreg_new<50> , \inreg_new<49> , \inreg_new<48> , \inreg_new<47> , \inreg_new<46> , \inreg_new<45> , \inreg_new<44> , \inreg_new<43> , \inreg_new<42> , \inreg_new<41> , \inreg_new<40> , \inreg_new<39> , \inreg_new<38> , \inreg_new<37> , \inreg_new<36> , \inreg_new<35> , \inreg_new<34> , \inreg_new<33> , \inreg_new<32> , \inreg_new<31> , \inreg_new<30> , \inreg_new<29> , \inreg_new<28> , \inreg_new<27> , \inreg_new<26> , \inreg_new<25> , \inreg_new<24> , \inreg_new<23> , \inreg_new<22> , \inreg_new<21> , \inreg_new<20> , \inreg_new<19> , \inreg_new<18> , \inreg_new<17> , \inreg_new<16> , \inreg_new<15> , \inreg_new<14> , \inreg_new<13> , \inreg_new<12> , \inreg_new<11> , \inreg_new<10> , \inreg_new<9> , \inreg_new<8> , \inreg_new<7> , \inreg_new<6> , \inreg_new<5> , \inreg_new<4> , \inreg_new<3> , \inreg_new<2> , \inreg_new<1> , \inreg_new<0> , \outreg_new<63> , \outreg_new<62> , \outreg_new<61> , \outreg_new<60> , \outreg_new<59> , \outreg_new<58> , \outreg_new<57> , \outreg_new<56> , \outreg_new<55> , \outreg_new<54> , \outreg_new<53> , \outreg_new<52> , \outreg_new<51> , \outreg_new<50> , \outreg_new<49> , \outreg_new<48> , \outreg_new<47> , \outreg_new<46> , \outreg_new<45> , \outreg_new<44> , \outreg_new<43> , \outreg_new<42> , \outreg_new<41> , \outreg_new<40> , \outreg_new<39> , \outreg_new<38> , \outreg_new<37> , \outreg_new<36> , \outreg_new<35> , \outreg_new<34> , \outreg_new<33> , \outreg_new<32> , \outreg_new<31> , \outreg_new<30> , \outreg_new<29> , \outreg_new<28> , \outreg_new<27> , \outreg_new<26> , \outreg_new<25> , \outreg_new<24> , \outreg_new<23> , \outreg_new<22> , \outreg_new<21> , \outreg_new<20> , \outreg_new<19> , \outreg_new<18> , \outreg_new<17> , \outreg_new<16> , \outreg_new<15> , \outreg_new<14> , \outreg_new<13> , \outreg_new<12> , \outreg_new<11> , \outreg_new<10> , \outreg_new<9> , \outreg_new<8> , \outreg_new<7> , \outreg_new<6> , \outreg_new<5> , \outreg_new<4> , \outreg_new<3> , \outreg_new<2> , \outreg_new<1> , \outreg_new<0> , \data_new<63> , \data_new<62> , \data_new<61> , \data_new<60> , \data_new<59> , \data_new<58> , \data_new<57> , \data_new<56> , \data_new<55> , \data_new<54> , \data_new<53> , \data_new<52> , \data_new<51> , \data_new<50> , \data_new<49> , \data_new<48> , \data_new<47> , \data_new<46> , \data_new<45> , \data_new<44> , \data_new<43> , \data_new<42> , \data_new<41> , \data_new<40> , \data_new<39> , \data_new<38> , \data_new<37> , \data_new<36> , \data_new<35> , \data_new<34> , \data_new<33> , \data_new<32> , \data_new<31> , \data_new<30> , \data_new<29> , \data_new<28> , \data_new<27> , \data_new<26> , \data_new<25> , \data_new<24> , \data_new<23> , \data_new<22> , \data_new<21> , \data_new<20> , \data_new<19> , \data_new<18> , \data_new<17> , \data_new<16> , \data_new<15> , \data_new<14> , \data_new<13> , \data_new<12> , \data_new<11> , \data_new<10> , \data_new<9> , \data_new<8> , \data_new<7> , \data_new<6> , \data_new<5> , \data_new<4> , \data_new<3> , \data_new<2> , \data_new<1> , \data_new<0> , \count_new<3> , \count_new<2> , \count_new<1> , \count_new<0> , \C_new<27> , \C_new<26> , \C_new<25> , \C_new<24> , \C_new<23> , \C_new<22> , \C_new<21> , \C_new<20> , \C_new<19> , \C_new<18> , \C_new<17> , \C_new<16> , \C_new<15> , \C_new<14> , \C_new<13> , \C_new<12> , \C_new<11> , \C_new<10> , \C_new<9> , \C_new<8> , \C_new<7> , \C_new<6> , \C_new<5> , \C_new<4> , \C_new<3> , \C_new<2> , \C_new<1> , \C_new<0> , \D_new<27> , \D_new<26> , \D_new<25> , \D_new<24> , \D_new<23> , \D_new<22> , \D_new<21> , \D_new<20> , \D_new<19> , \D_new<18> , \D_new<17> , \D_new<16> , \D_new<15> , \D_new<14> , \D_new<13> , \D_new<12> , \D_new<11> , \D_new<10> , \D_new<9> , \D_new<8> , \D_new<7> , \D_new<6> , \D_new<5> , \D_new<4> , \D_new<3> , \D_new<2> , \D_new<1> , \D_new<0> , \encrypt_mode_new<0> );
input
  \data<63> ,
  \data<61> ,
  \data<62> ,
  \reset<0> ,
  \outreg<58> ,
  \inreg<0> ,
  \outreg<57> ,
  \inreg<1> ,
  \outreg<56> ,
  \inreg<2> ,
  \outreg<55> ,
  \inreg<3> ,
  \inreg<4> ,
  \inreg<5> ,
  \inreg<6> ,
  \outreg<59> ,
  \inreg<7> ,
  \outreg<50> ,
  \inreg<8> ,
  \inreg<9> ,
  \outreg<54> ,
  \outreg<53> ,
  \outreg<52> ,
  \outreg<51> ,
  \load_key<0> ,
  \outreg<60> ,
  \outreg<63> ,
  \outreg<62> ,
  \outreg<61> ,
  \D<0> ,
  \D<1> ,
  \D<2> ,
  \D<3> ,
  \D<4> ,
  \D<5> ,
  \D<6> ,
  \C<10> ,
  \D<7> ,
  \C<11> ,
  \D<8> ,
  \C<12> ,
  \D<9> ,
  \C<13> ,
  \C<14> ,
  \C<15> ,
  \C<16> ,
  \C<17> ,
  \C<18> ,
  \C<19> ,
  \outreg<18> ,
  \outreg<17> ,
  \outreg<16> ,
  \outreg<15> ,
  \C<20> ,
  \outreg<19> ,
  \C<21> ,
  \outreg<10> ,
  \C<22> ,
  \C<23> ,
  \C<24> ,
  \C<25> ,
  \outreg<14> ,
  \C<26> ,
  \outreg<13> ,
  \C<27> ,
  \outreg<12> ,
  \outreg<11> ,
  \outreg<28> ,
  \outreg<27> ,
  \outreg<26> ,
  \outreg<25> ,
  \outreg<29> ,
  \outreg<20> ,
  \data<3> ,
  \data<4> ,
  \data<1> ,
  \outreg<24> ,
  \data<2> ,
  \outreg<23> ,
  \outreg<22> ,
  \data<0> ,
  \outreg<21> ,
  \outreg<38> ,
  \outreg<37> ,
  \outreg<36> ,
  \outreg<35> ,
  \data<9> ,
  \data<7> ,
  \data<8> ,
  \outreg<39> ,
  \data<5> ,
  \outreg<30> ,
  \data<6> ,
  \outreg<34> ,
  \outreg<33> ,
  \outreg<32> ,
  \outreg<31> ,
  \outreg<48> ,
  \outreg<47> ,
  \outreg<46> ,
  \outreg<45> ,
  \outreg<49> ,
  \outreg<40> ,
  \outreg<44> ,
  \outreg<43> ,
  \outreg<42> ,
  \outreg<41> ,
  \D<10> ,
  \D<11> ,
  \D<12> ,
  \D<13> ,
  \D<14> ,
  \D<15> ,
  \D<16> ,
  \D<17> ,
  \D<18> ,
  \D<19> ,
  \D<20> ,
  \D<21> ,
  \data_in<7> ,
  \D<22> ,
  \D<23> ,
  \data_in<5> ,
  \D<24> ,
  \data_in<6> ,
  \D<25> ,
  \D<26> ,
  \D<27> ,
  \data_in<0> ,
  \data_in<3> ,
  \data_in<4> ,
  \data_in<1> ,
  \data_in<2> ,
  \data<37> ,
  \data<38> ,
  \data<35> ,
  \data<36> ,
  \data<39> ,
  \data<30> ,
  \data<33> ,
  \data<34> ,
  \data<31> ,
  \data<32> ,
  \data<47> ,
  \data<48> ,
  \data<45> ,
  \data<46> ,
  \data<49> ,
  \data<40> ,
  \data<43> ,
  \data<44> ,
  \data<41> ,
  \data<42> ,
  \data<17> ,
  \data<18> ,
  \data<15> ,
  \count<0> ,
  \data<16> ,
  \count<3> ,
  \data<19> ,
  \count<1> ,
  \count<2> ,
  \data<10> ,
  \data<13> ,
  \data<14> ,
  \data<11> ,
  \data<12> ,
  \data<27> ,
  \data<28> ,
  \data<25> ,
  \data<26> ,
  \data<29> ,
  \data<20> ,
  \data<23> ,
  \data<24> ,
  \data<21> ,
  \data<22> ,
  \C<0> ,
  \C<1> ,
  \C<2> ,
  \C<3> ,
  \C<4> ,
  \C<5> ,
  \C<6> ,
  \C<7> ,
  \C<8> ,
  \C<9> ,
  \inreg<12> ,
  \inreg<11> ,
  \inreg<14> ,
  \inreg<13> ,
  \inreg<10> ,
  \inreg<19> ,
  \inreg<16> ,
  \inreg<15> ,
  \inreg<18> ,
  \inreg<17> ,
  \inreg<22> ,
  \inreg<21> ,
  \inreg<24> ,
  \inreg<23> ,
  \inreg<20> ,
  \inreg<29> ,
  \inreg<26> ,
  \inreg<25> ,
  \outreg<9> ,
  \inreg<28> ,
  \inreg<27> ,
  \inreg<32> ,
  \inreg<31> ,
  \outreg<5> ,
  \inreg<34> ,
  \outreg<6> ,
  \inreg<33> ,
  \outreg<7> ,
  \outreg<8> ,
  \outreg<1> ,
  \inreg<30> ,
  \outreg<2> ,
  \outreg<3> ,
  \outreg<4> ,
  \inreg<39> ,
  \inreg<36> ,
  \outreg<0> ,
  \inreg<35> ,
  \inreg<38> ,
  \inreg<37> ,
  \inreg<42> ,
  \inreg<41> ,
  \inreg<44> ,
  \inreg<43> ,
  \inreg<40> ,
  \inreg<49> ,
  \inreg<46> ,
  \inreg<45> ,
  \encrypt_mode<0> ,
  \inreg<48> ,
  \inreg<47> ,
  \inreg<52> ,
  \inreg<51> ,
  \inreg<54> ,
  \inreg<53> ,
  \inreg<50> ,
  \inreg<55> ,
  \data<57> ,
  \data<58> ,
  \data<55> ,
  \data<56> ,
  \encrypt<0> ,
  \data<59> ,
  \data<50> ,
  \data<53> ,
  \data<54> ,
  \data<51> ,
  \data<52> ,
  \data<60> ;
output
  \data_new<25> ,
  \inreg_new<45> ,
  \data_new<26> ,
  \data_new<13> ,
  \data_new<14> ,
  \data_new<11> ,
  \inreg_new<49> ,
  \data_new<12> ,
  \inreg_new<30> ,
  \outreg_new<11> ,
  \count_new<0> ,
  \outreg_new<12> ,
  \data_new<10> ,
  \outreg_new<13> ,
  \outreg_new<14> ,
  \inreg_new<34> ,
  \count_new<3> ,
  \inreg_new<33> ,
  \inreg_new<32> ,
  \count_new<1> ,
  \data_new<19> ,
  \inreg_new<31> ,
  \count_new<2> ,
  \outreg_new<10> ,
  \inreg_new<38> ,
  \outreg_new<19> ,
  \data_new<17> ,
  \inreg_new<37> ,
  \data_new<18> ,
  \inreg_new<36> ,
  \data_new<15> ,
  \inreg_new<35> ,
  \data_new<16> ,
  \outreg_new<15> ,
  \outreg_new<16> ,
  \outreg_new<17> ,
  \inreg_new<39> ,
  \outreg_new<18> ,
  \outreg_new<21> ,
  \outreg_new<22> ,
  \outreg_new<23> ,
  \outreg_new<24> ,
  \outreg_new<20> ,
  \outreg_new<29> ,
  \outreg_new<25> ,
  \outreg_new<26> ,
  \outreg_new<27> ,
  \outreg_new<28> ,
  \outreg_new<31> ,
  \outreg_new<32> ,
  \outreg_new<33> ,
  \outreg_new<34> ,
  \outreg_new<30> ,
  \outreg_new<39> ,
  \outreg_new<35> ,
  \outreg_new<36> ,
  \outreg_new<37> ,
  \outreg_new<38> ,
  \outreg_new<41> ,
  \outreg_new<42> ,
  \outreg_new<43> ,
  \outreg_new<44> ,
  \outreg_new<40> ,
  \outreg_new<49> ,
  \outreg_new<45> ,
  \outreg_new<46> ,
  \outreg_new<47> ,
  \outreg_new<48> ,
  \C_new<23> ,
  \C_new<24> ,
  \C_new<21> ,
  \C_new<22> ,
  \C_new<20> ,
  \data_new<4> ,
  \data_new<3> ,
  \C_new<27> ,
  \data_new<2> ,
  \data_new<1> ,
  \C_new<25> ,
  \data_new<0> ,
  \C_new<26> ,
  \C_new<13> ,
  \C_new<14> ,
  \C_new<11> ,
  \C_new<12> ,
  \C_new<10> ,
  \data_new<9> ,
  \data_new<8> ,
  \data_new<7> ,
  \data_new<6> ,
  \data_new<5> ,
  \C_new<19> ,
  \C_new<17> ,
  \C_new<18> ,
  \C_new<15> ,
  \C_new<16> ,
  \D_new<13> ,
  \D_new<14> ,
  \D_new<11> ,
  \D_new<12> ,
  \D_new<10> ,
  \data_new<63> ,
  \data_new<61> ,
  \data_new<62> ,
  \D_new<19> ,
  \data_new<60> ,
  \D_new<17> ,
  \D_new<18> ,
  \D_new<15> ,
  \D_new<16> ,
  \D_new<23> ,
  \D_new<24> ,
  \D_new<21> ,
  \D_new<22> ,
  \D_new<20> ,
  \data_new<53> ,
  \data_new<54> ,
  \data_new<51> ,
  \data_new<52> ,
  \data_new<50> ,
  \D_new<27> ,
  \D_new<25> ,
  \D_new<26> ,
  \data_new<59> ,
  \data_new<57> ,
  \data_new<58> ,
  \data_new<55> ,
  \data_new<56> ,
  \D_new<7> ,
  \C_new<6> ,
  \D_new<8> ,
  \C_new<5> ,
  \D_new<5> ,
  \C_new<8> ,
  \D_new<6> ,
  \C_new<7> ,
  \C_new<9> ,
  \D_new<9> ,
  \D_new<0> ,
  \C_new<0> ,
  \D_new<3> ,
  \C_new<2> ,
  \D_new<4> ,
  \C_new<1> ,
  \D_new<1> ,
  \C_new<4> ,
  \D_new<2> ,
  \C_new<3> ,
  \inreg_new<50> ,
  \inreg_new<9> ,
  \inreg_new<54> ,
  \inreg_new<53> ,
  \inreg_new<52> ,
  \inreg_new<6> ,
  \inreg_new<51> ,
  \inreg_new<5> ,
  \inreg_new<8> ,
  \inreg_new<7> ,
  \inreg_new<2> ,
  \inreg_new<55> ,
  \inreg_new<1> ,
  \inreg_new<4> ,
  \inreg_new<3> ,
  \inreg_new<0> ,
  \encrypt_mode_new<0> ,
  \outreg_new<9> ,
  \outreg_new<51> ,
  \outreg_new<52> ,
  \outreg_new<53> ,
  \outreg_new<5> ,
  \outreg_new<54> ,
  \outreg_new<6> ,
  \outreg_new<7> ,
  \outreg_new<8> ,
  \outreg_new<1> ,
  \outreg_new<50> ,
  \outreg_new<2> ,
  \outreg_new<59> ,
  \outreg_new<3> ,
  \outreg_new<4> ,
  \outreg_new<55> ,
  \data_new<43> ,
  \outreg_new<56> ,
  \data_new<44> ,
  \outreg_new<0> ,
  \outreg_new<57> ,
  \data_new<41> ,
  \outreg_new<58> ,
  \data_new<42> ,
  \inreg_new<20> ,
  \outreg_new<61> ,
  \outreg_new<62> ,
  \data_new<40> ,
  \outreg_new<63> ,
  \inreg_new<24> ,
  \inreg_new<23> ,
  \inreg_new<22> ,
  \data_new<49> ,
  \inreg_new<21> ,
  \outreg_new<60> ,
  \inreg_new<28> ,
  \data_new<47> ,
  \inreg_new<27> ,
  \data_new<48> ,
  \inreg_new<26> ,
  \data_new<45> ,
  \inreg_new<25> ,
  \data_new<46> ,
  \data_new<33> ,
  \data_new<34> ,
  \data_new<31> ,
  \inreg_new<29> ,
  \data_new<32> ,
  \inreg_new<10> ,
  \data_new<30> ,
  \inreg_new<14> ,
  \inreg_new<13> ,
  \inreg_new<12> ,
  \data_new<39> ,
  \inreg_new<11> ,
  \inreg_new<18> ,
  \data_new<37> ,
  \inreg_new<17> ,
  \data_new<38> ,
  \inreg_new<16> ,
  \data_new<35> ,
  \inreg_new<15> ,
  \data_new<36> ,
  \data_new<23> ,
  \data_new<24> ,
  \data_new<21> ,
  \inreg_new<19> ,
  \data_new<22> ,
  \inreg_new<40> ,
  \data_new<20> ,
  \inreg_new<44> ,
  \inreg_new<43> ,
  \inreg_new<42> ,
  \data_new<29> ,
  \inreg_new<41> ,
  \inreg_new<48> ,
  \data_new<27> ,
  \inreg_new<47> ,
  \data_new<28> ,
  \inreg_new<46> ;
wire
  \$$COND258<0>226.1 ,
  \[568] ,
  \$$COND216<0>226.1 ,
  \$$COND365<0>376.1 ,
  \$$COND180<0>151.1 ,
  \[189] ,
  \[569] ,
  \$$COND391<0>451.1 ,
  \[190] ,
  \[570] ,
  \[191] ,
  \[571] ,
  \[192] ,
  \[572] ,
  \[193] ,
  \main_1/preS<28>0.1 ,
  \[573] ,
  \[194] ,
  \[574] ,
  \[195] ,
  \[575] ,
  \main_1/S7_1/$S7<3>526.1 ,
  \[196] ,
  \[576] ,
  \main_1/preS<11>0.1 ,
  \[197] ,
  \[577] ,
  \[198] ,
  \[578] ,
  \$$COND328<0>376.1 ,
  \[199] ,
  \[579] ,
  \$$COND521<0>601.1 ,
  \main_1/preS<7>0.1 ,
  \[1] ,
  \[580] ,
  \[2] ,
  \[581] ,
  \[3] ,
  \[582] ,
  \[4] ,
  \[583] ,
  \main_1/S2_1/$S2<1>151.1 ,
  \[5] ,
  \[584] ,
  \[6] ,
  \[585] ,
  \[7] ,
  \[586] ,
  \[8] ,
  \[587] ,
  \[9] ,
  \[588] ,
  \[589] ,
  \main_1/preS<24>0.1 ,
  \main_1/S0_1/$S0<2>1.1 ,
  \main_1/S3_1/$S3<3>226.1 ,
  \main_1/S4_1/$S4<2>301.1 ,
  \main_1/S1_1/$S1<3>76.1 ,
  \$$COND34<0>1.1 ,
  \[590] ,
  \main_1/preS<36>0.1 ,
  \[591] ,
  \[592] ,
  \[593] ,
  \[594] ,
  \[595] ,
  \[596] ,
  \[597] ,
  \[598] ,
  \$$COND238<0>226.1 ,
  \[599] ,
  \$$COND95<0>76.1 ,
  \main_1/preS<20>0.1 ,
  \$$COND99<0>76.1 ,
  \main_1/preS<2>0.1 ,
  \main_1/preS<32>0.1 ,
  \$$COND196<0>226.1 ,
  \main_1/S5_1/$S5<0>376.1 ,
  \main_1/preS<45>0.1 ,
  \$$COND76<0>76.1 ,
  \$$COND484<0>526.1 ,
  \$$COND70<0>76.1 ,
  \main_1/preS<18>0.1 ,
  \main_1/preS<41>0.1 ,
  \main_1/S4_1/$S4<1>301.1 ,
  \$$COND43<0>1.1 ,
  \main_1/S6_1/$S6<0>451.1 ,
  \$$COND82<0>76.1 ,
  \$$COND157<0>151.1 ,
  \$$COND307<0>301.1 ,
  \[200] ,
  \[201] ,
  \[202] ,
  \main_1/preS<14>0.1 ,
  \[203] ,
  \[204] ,
  \[205] ,
  \[206] ,
  \main_1/preS<6>0.1 ,
  \[207] ,
  \[208] ,
  \[209] ,
  \$$COND65<0>76.1 ,
  \[210] ,
  \[211] ,
  \[212] ,
  \[213] ,
  \[214] ,
  \main_1/preS<27>0.1 ,
  \[215] ,
  \[216] ,
  \$$COND281<0>301.1 ,
  \[217] ,
  \main_1/S0_1/$S0<3>1.1 ,
  \[218] ,
  \main_1/preS<10>0.1 ,
  \[219] ,
  \$$COND311<0>301.1 ,
  \main_1/preS<39>0.1 ,
  \[220] ,
  \[600] ,
  \[221] ,
  \[601] ,
  \[222] ,
  \[602] ,
  \[223] ,
  \[603] ,
  \[224] ,
  \[604] ,
  \[225] ,
  \[605] ,
  \[226] ,
  \[606] ,
  \[227] ,
  \[607] ,
  \[228] ,
  \[608] ,
  \$$COND371<0>376.1 ,
  \[229] ,
  \[609] ,
  \main_1/S2_1/$S2<3>151.1 ,
  \main_1/preS<23>0.1 ,
  \main_1/S5_1/$S5<2>376.1 ,
  \[230] ,
  \[610] ,
  \[231] ,
  \[611] ,
  \[232] ,
  \main_1/preS<35>0.1 ,
  \[612] ,
  \[233] ,
  \[613] ,
  \[234] ,
  \[614] ,
  \[235] ,
  \[615] ,
  \[236] ,
  \[616] ,
  \[237] ,
  \[617] ,
  \[238] ,
  \[618] ,
  \[239] ,
  \[619] ,
  \[240] ,
  \[620] ,
  \[241] ,
  \[621] ,
  \[242] ,
  \[622] ,
  \[243] ,
  \[623] ,
  \[244] ,
  \[624] ,
  \[245] ,
  \[625] ,
  \main_1/preS<1>0.1 ,
  \[626] ,
  \[627] ,
  \[628] ,
  \main_1/preS<31>0.1 ,
  \[629] ,
  \main_1/S6_1/$S6<2>451.1 ,
  \[630] ,
  \[631] ,
  \[632] ,
  \[633] ,
  \[634] ,
  \[635] ,
  \[636] ,
  \[637] ,
  \[638] ,
  \[639] ,
  \main_1/preS<44>0.1 ,
  \main_1/S7_1/$S7<0>526.1 ,
  \[640] ,
  \main_1/S1_1/$S1<1>76.1 ,
  \[641] ,
  \[642] ,
  \[643] ,
  \[644] ,
  \[645] ,
  \[646] ,
  \[647] ,
  \[648] ,
  \$$COND225<0>226.1 ,
  \$$COND354<0>376.1 ,
  \$$COND244<0>226.1 ,
  \[649] ,
  \main_1/preS<17>0.1 ,
  \[650] ,
  \main_1/S5_1/$S5<1>376.1 ,
  \main_1/preS<40>0.1 ,
  \[651] ,
  \main_1/preS<9>0.1 ,
  \[652] ,
  \[653] ,
  \[654] ,
  \[655] ,
  \[656] ,
  \[657] ,
  \main_1/S3_1/$S3<0>226.1 ,
  \main_1/S4_1/$S4<3>301.1 ,
  \[658] ,
  \[659] ,
  \[660] ,
  \[661] ,
  \$$COND520<0>0.1 ,
  \[662] ,
  \main_1/S0_1/$S0<0>1.1 ,
  \[663] ,
  \main_1/preS<13>0.1 ,
  \[664] ,
  \[665] ,
  \[666] ,
  \[667] ,
  \$$COND414<0>451.1 ,
  \main_1/preS<5>0.1 ,
  \[668] ,
  \[669] ,
  \[670] ,
  \[671] ,
  \main_1/S6_1/$S6<1>451.1 ,
  \[672] ,
  \[673] ,
  \[674] ,
  \main_1/S1_1/$S1<0>76.1 ,
  \[675] ,
  \main_1/preS<26>0.1 ,
  \[676] ,
  \[677] ,
  \[678] ,
  \[679] ,
  \main_1/preS<38>0.1 ,
  \[490] ,
  \[491] ,
  \[492] ,
  \[682] ,
  \[493] ,
  \[494] ,
  \[495] ,
  \[496] ,
  \[497] ,
  \[498] ,
  \$$COND358<0>376.1 ,
  \[499] ,
  \main_1/preS<22>0.1 ,
  \generate_key_1/freeze<0>605.1 ,
  \[693] ,
  \main_1/preS<34>0.1 ,
  \$$COND359<0>376.1 ,
  \$$COND249<0>226.1 ,
  \$$COND207<0>226.1 ,
  \main_1/S1_1/$S1<2>76.1 ,
  \main_1/S7_1/$S7<2>526.1 ,
  \$$COND40<0>1.1 ,
  \main_1/preS<47>0.1 ,
  \main_1/preS<4>0.1 ,
  \main_1/preS<30>0.1 ,
  \main_1/S3_1/$S3<2>226.1 ,
  \[10] ,
  \[11] ,
  \[12] ,
  \[13] ,
  \[14] ,
  \[15] ,
  \main_1/preS<43>0.1 ,
  \[16] ,
  \main_1/preS<0>0.1 ,
  \[17] ,
  \[18] ,
  \[19] ,
  \[20] ,
  \[21] ,
  \[22] ,
  \[23] ,
  \[24] ,
  \[25] ,
  \[26] ,
  \[27] ,
  \[28] ,
  \main_1/preS<16>0.1 ,
  \[100] ,
  \[29] ,
  \[101] ,
  \[102] ,
  \[103] ,
  \[104] ,
  \main_1/S2_1/$S2<0>151.1 ,
  \[105] ,
  \[106] ,
  \[107] ,
  \[30] ,
  \main_1/S5_1/$S5<3>376.1 ,
  \[108] ,
  \[31] ,
  \[109] ,
  \[32] ,
  \[33] ,
  \[34] ,
  \[35] ,
  \[36] ,
  \[37] ,
  \main_1/S7_1/$S7<1>526.1 ,
  \[38] ,
  \[110] ,
  \[39] ,
  \[111] ,
  \main_1/preS<29>0.1 ,
  \[112] ,
  \[113] ,
  \[114] ,
  \[115] ,
  \main_1/preS<12>0.1 ,
  \[116] ,
  \[117] ,
  \[40] ,
  \[118] ,
  \[41] ,
  \$$COND445<0>451.1 ,
  \[119] ,
  \[42] ,
  \main_1/preS<8>0.1 ,
  \[43] ,
  \[44] ,
  \[45] ,
  \[46] ,
  \$$COND477<0>526.1 ,
  \[47] ,
  \[48] ,
  \[120] ,
  \[49] ,
  \[500] ,
  \[121] ,
  \[501] ,
  \[122] ,
  \[502] ,
  \[123] ,
  \[503] ,
  \[124] ,
  \[504] ,
  \[125] ,
  \[505] ,
  \[126] ,
  \main_1/S3_1/$S3<1>226.1 ,
  \[506] ,
  \[127] ,
  \[50] ,
  \[507] ,
  \main_1/preS<25>0.1 ,
  \[128] ,
  \[51] ,
  \[508] ,
  \$$COND210<0>226.1 ,
  \main_1/S6_1/$S6<3>451.1 ,
  \[129] ,
  \[52] ,
  \[509] ,
  \[53] ,
  \main_1/S0_1/$S0<1>1.1 ,
  \[54] ,
  \[55] ,
  \[56] ,
  \[57] ,
  \[58] ,
  \main_1/preS<37>0.1 ,
  \[130] ,
  \[59] ,
  \[510] ,
  \[131] ,
  \[511] ,
  \[701] ,
  \[132] ,
  \[512] ,
  \[702] ,
  \[133] ,
  \[513] ,
  \[703] ,
  \[134] ,
  \[514] ,
  \[704] ,
  \[135] ,
  \[515] ,
  \[705] ,
  \[136] ,
  \[516] ,
  \[706] ,
  \[137] ,
  \[60] ,
  \[517] ,
  \[707] ,
  \[138] ,
  \[61] ,
  \[518] ,
  \[139] ,
  \[62] ,
  \$$COND317<0>301.1 ,
  \[519] ,
  \[709] ,
  \[63] ,
  \[64] ,
  \[65] ,
  \[66] ,
  \[67] ,
  \main_1/preS<21>0.1 ,
  \[68] ,
  \[140] ,
  \[69] ,
  \[520] ,
  \[710] ,
  \[141] ,
  \generate_key_1/shift_by_one<0>605.1 ,
  \[521] ,
  \[711] ,
  \[142] ,
  \[522] ,
  \[712] ,
  \[143] ,
  \[523] ,
  \[713] ,
  \[144] ,
  \[524] ,
  \[714] ,
  \[145] ,
  \[525] ,
  \main_1/preS<33>0.1 ,
  \[715] ,
  \[146] ,
  \$$COND286<0>301.1 ,
  \[526] ,
  \[716] ,
  \[147] ,
  \[70] ,
  \[527] ,
  \[717] ,
  \[148] ,
  \[71] ,
  \$$COND254<0>226.1 ,
  \[528] ,
  \[718] ,
  \[149] ,
  \[72] ,
  \[529] ,
  \[719] ,
  \[73] ,
  \[74] ,
  \[75] ,
  \[76] ,
  \[77] ,
  \[78] ,
  \[150] ,
  \[79] ,
  \[530] ,
  \[720] ,
  \[151] ,
  \[531] ,
  \[721] ,
  \[152] ,
  \[532] ,
  \[722] ,
  \main_1/S4_1/$S4<0>301.1 ,
  \[153] ,
  \[533] ,
  \[723] ,
  \[154] ,
  \[534] ,
  \[724] ,
  \[155] ,
  \[535] ,
  \[725] ,
  \[156] ,
  \[536] ,
  \[726] ,
  \[157] ,
  \[80] ,
  \[537] ,
  \[727] ,
  \main_1/preS<46>0.1 ,
  \[158] ,
  \[81] ,
  \[538] ,
  \[728] ,
  \$$COND232<0>226.1 ,
  \main_1/preS<3>0.1 ,
  \[159] ,
  \[82] ,
  \[539] ,
  \[729] ,
  \[83] ,
  \[84] ,
  \[85] ,
  \[86] ,
  \[87] ,
  \[88] ,
  \[160] ,
  \main_1/S2_1/$S2<2>151.1 ,
  \[89] ,
  \[540] ,
  \[730] ,
  \[161] ,
  \[541] ,
  \[731] ,
  \[162] ,
  \[542] ,
  \[732] ,
  \[163] ,
  \[543] ,
  \[164] ,
  \[544] ,
  \[165] ,
  \[545] ,
  \[166] ,
  \[546] ,
  \[167] ,
  \[90] ,
  \[547] ,
  \[168] ,
  \[91] ,
  \[548] ,
  \$$COND233<0>226.1 ,
  \[169] ,
  \[92] ,
  \[549] ,
  \[93] ,
  \main_1/preS<19>0.1 ,
  \[94] ,
  \[95] ,
  \[96] ,
  \[97] ,
  \main_1/preS<42>0.1 ,
  \[98] ,
  \[170] ,
  \[99] ,
  \[550] ,
  \[171] ,
  \[551] ,
  \[172] ,
  \[552] ,
  \[173] ,
  \[553] ,
  \[174] ,
  \[554] ,
  \[175] ,
  \[555] ,
  \[176] ,
  \[556] ,
  \[177] ,
  \[557] ,
  \[178] ,
  \[558] ,
  \[179] ,
  \[559] ,
  \[180] ,
  \[560] ,
  \main_1/preS<15>0.1 ,
  \[181] ,
  \[561] ,
  \[182] ,
  \[562] ,
  \[183] ,
  \[184] ,
  \[564] ,
  \[185] ,
  \[565] ,
  \[186] ,
  \[566] ,
  \[187] ,
  \[567] ,
  \[188] ;
assign
  \$$COND258<0>226.1  = \[551]  & (\[529]  & ~\[510] ),
  \[568]  = ~\main_1/preS<8>0.1  & ~\main_1/preS<6>0.1 ,
  \data_new<25>  = \[159] ,
  \$$COND216<0>226.1  = \[729]  & \[712] ,
  \inreg_new<45>  = \[11] ,
  \$$COND365<0>376.1  = \[635]  & (\[531]  & ~\main_1/preS<32>0.1 ),
  \$$COND180<0>151.1  = \[715]  & \[656] ,
  \[189]  = (\[503]  & \C<26> ) | ((\[502]  & \C<0> ) | ((\[501]  & \C<1> ) | ((\[500]  & \C<25> ) | ((\[499]  & \C<27> ) | ((\[498]  & \inreg<48> ) | (\[497]  & \inreg<27> )))))),
  \[569]  = \[531]  & \main_1/preS<35>0.1 ,
  \data_new<26>  = \[158] ,
  \data_new<13>  = \[171] ,
  \$$COND391<0>451.1  = \[727]  & \[638] ,
  \data_new<14>  = \[170] ,
  \data_new<11>  = \[173] ,
  \inreg_new<49>  = \[7] ,
  \data_new<12>  = \[172] ,
  \inreg_new<30>  = \[26] ,
  \outreg_new<11>  = \[109] ,
  \count_new<0>  = \[188] ,
  \outreg_new<12>  = \[108] ,
  \data_new<10>  = \[174] ,
  \[190]  = (\[503]  & \C<25> ) | ((\[502]  & \C<27> ) | ((\[501]  & \C<0> ) | ((\[500]  & \C<24> ) | ((\[499]  & \C<26> ) | ((\[498]  & \inreg<27> ) | (\[497]  & \inreg<35> )))))),
  \outreg_new<13>  = \[107] ,
  \[570]  = ~\[515]  & ~\main_1/preS<10>0.1 ,
  \[191]  = (\[503]  & \C<24> ) | ((\[502]  & \C<26> ) | ((\[501]  & \C<27> ) | ((\[500]  & \C<23> ) | ((\[499]  & \C<25> ) | ((\[498]  & \inreg<35> ) | (\[497]  & \inreg<43> )))))),
  \outreg_new<14>  = \[106] ,
  \[571]  = \main_1/preS<8>0.1  & \main_1/preS<11>0.1 ,
  \inreg_new<34>  = \[22] ,
  \[192]  = (\[503]  & \C<23> ) | ((\[502]  & \C<25> ) | ((\[501]  & \C<26> ) | ((\[500]  & \C<22> ) | ((\[499]  & \C<24> ) | ((\[498]  & \inreg<43> ) | (\[497]  & \inreg<51> )))))),
  \count_new<3>  = \[185] ,
  \[572]  = \[529]  & ~\main_1/preS<21>0.1 ,
  \inreg_new<33>  = \[23] ,
  \[193]  = (\[503]  & \C<22> ) | ((\[502]  & \C<24> ) | ((\[501]  & \C<25> ) | ((\[500]  & \C<21> ) | ((\[499]  & \C<23> ) | ((\[498]  & \inreg<51> ) | (\[497]  & \data_in<2> )))))),
  \main_1/preS<28>0.1  = (~\data<51>  & \D<18> ) | (\data<51>  & ~\D<18> ),
  \[573]  = \main_1/preS<38>0.1  & ~\main_1/preS<37>0.1 ,
  \inreg_new<32>  = \[24] ,
  \[194]  = (\[503]  & \C<21> ) | ((\[502]  & \C<23> ) | ((\[501]  & \C<24> ) | ((\[500]  & \C<20> ) | ((\[499]  & \C<22> ) | ((\[498]  & \data_in<2> ) | (\[497]  & \inreg<2> )))))),
  \count_new<1>  = \[187] ,
  \[574]  = \main_1/preS<41>0.1  & ~\main_1/preS<40>0.1 ,
  \data_new<19>  = \[165] ,
  \inreg_new<31>  = \[25] ,
  \[195]  = (\[503]  & \C<20> ) | ((\[502]  & \C<22> ) | ((\[501]  & \C<23> ) | ((\[500]  & \C<19> ) | ((\[499]  & \C<21> ) | ((\[498]  & \inreg<2> ) | (\[497]  & \inreg<10> )))))),
  \count_new<2>  = \[186] ,
  \outreg_new<10>  = \[110] ,
  \[575]  = ~\main_1/preS<28>0.1  & \main_1/preS<24>0.1 ,
  \main_1/S7_1/$S7<3>526.1  = (~\[711]  & (~\[655]  & (\[580]  & (~\[564]  & ~\main_1/preS<42>0.1 )))) | ((~\[665]  & (~\[655]  & (~\[513]  & (~\main_1/preS<47>0.1  & \main_1/preS<42>0.1 )))) | ((~\[580]  & (\[564]  & (~\[549]  & (~\[517]  & ~\main_1/preS<45>0.1 )))) | ((~\[655]  & (\[583]  & (~\[564]  & \main_1/preS<43>0.1 ))) | ((\[655]  & (~\[583]  & (~\main_1/preS<47>0.1  & ~\main_1/preS<42>0.1 ))) | ((\[583]  & (~\main_1/preS<46>0.1  & (~\main_1/preS<43>0.1  & ~\$$COND477<0>526.1 ))) | ((~\[534]  & (\[513]  & (\main_1/preS<46>0.1  & \main_1/preS<43>0.1 ))) | ((\[534]  & (\[517]  & (~\main_1/preS<45>0.1  & \main_1/preS<43>0.1 ))) | ((\[665]  & (\[649]  & ~\main_1/preS<44>0.1 )) | ((\[655]  & (\[513]  & \main_1/preS<43>0.1 )) | ((\[580]  & (\[564]  & \main_1/preS<42>0.1 )) | ((\[580]  & (\[513]  & ~\main_1/preS<46>0.1 )) | (\[560]  & (\[513]  & ~\[511] ))))))))))))),
  \inreg_new<38>  = \[18] ,
  \[196]  = (\[503]  & \C<19> ) | ((\[502]  & \C<21> ) | ((\[501]  & \C<22> ) | ((\[500]  & \C<18> ) | ((\[499]  & \C<20> ) | ((\[498]  & \inreg<10> ) | (\[497]  & \inreg<18> )))))),
  \outreg_new<19>  = \[101] ,
  \[576]  = ~\main_1/preS<26>0.1  & \main_1/preS<25>0.1 ,
  \data_new<17>  = \[167] ,
  \inreg_new<37>  = \[19] ,
  \main_1/preS<11>0.1  = (~\data<40>  & \C<9> ) | (\data<40>  & ~\C<9> ),
  \[197]  = (\[503]  & \C<18> ) | ((\[502]  & \C<20> ) | ((\[501]  & \C<21> ) | ((\[500]  & \C<17> ) | ((\[499]  & \C<19> ) | ((\[498]  & \inreg<18> ) | (\[497]  & \inreg<26> )))))),
  \[577]  = \main_1/preS<40>0.1  & \main_1/preS<39>0.1 ,
  \data_new<18>  = \[166] ,
  \inreg_new<36>  = \[20] ,
  \[198]  = (\[503]  & \C<17> ) | ((\[502]  & \C<19> ) | ((\[501]  & \C<20> ) | ((\[500]  & \C<16> ) | ((\[499]  & \C<18> ) | ((\[498]  & \inreg<26> ) | (\[497]  & \inreg<34> )))))),
  \[578]  = ~\main_1/preS<34>0.1  & \main_1/preS<33>0.1 ,
  \data_new<15>  = \[169] ,
  \$$COND328<0>376.1  = \[701]  & ~\[505] ,
  \inreg_new<35>  = \[21] ,
  \[199]  = (\[503]  & \C<16> ) | ((\[502]  & \C<18> ) | ((\[501]  & \C<19> ) | ((\[500]  & \C<15> ) | ((\[499]  & \C<17> ) | ((\[498]  & \inreg<34> ) | (\[497]  & \inreg<42> )))))),
  \[579]  = ~\[510]  & ~\main_1/preS<20>0.1 ,
  \data_new<16>  = \[168] ,
  \outreg_new<15>  = \[105] ,
  \$$COND521<0>601.1  = \$$COND520<0>0.1  & \load_key<0> ,
  \outreg_new<16>  = \[104] ,
  \main_1/preS<7>0.1  = (~\data<36>  & \C<27> ) | (\data<36>  & ~\C<27> ),
  \outreg_new<17>  = \[103] ,
  \inreg_new<39>  = \[17] ,
  \outreg_new<18>  = \[102] ,
  \outreg_new<21>  = \[99] ,
  \outreg_new<22>  = \[98] ,
  \[1]  = (\[493]  & \inreg<47> ) | (\[492]  & \inreg<55> ),
  \outreg_new<23>  = \[97] ,
  \[580]  = \main_1/preS<47>0.1  & ~\main_1/preS<43>0.1 ,
  \[2]  = (\[493]  & \inreg<46> ) | (\[492]  & \inreg<54> ),
  \outreg_new<24>  = \[96] ,
  \[581]  = ~\main_1/preS<26>0.1  & ~\main_1/preS<25>0.1 ,
  \[3]  = (\[493]  & \inreg<45> ) | (\[492]  & \inreg<53> ),
  \[582]  = \main_1/preS<15>0.1  & \main_1/preS<13>0.1 ,
  \[4]  = (\[493]  & \inreg<44> ) | (\[492]  & \inreg<52> ),
  \[583]  = \main_1/preS<45>0.1  & ~\main_1/preS<42>0.1 ,
  \main_1/S2_1/$S2<1>151.1  = (~\[715]  & (~\[672]  & (~\[617]  & (~\[555]  & (~\main_1/preS<15>0.1  & ~\main_1/preS<14>0.1 ))))) | ((\[676]  & (~\[541]  & (~\[530]  & \[519] ))) | ((\[676]  & (\[672]  & ~\[519] )) | ((\[676]  & (\[530]  & \main_1/preS<16>0.1 )) | ((\[623]  & (\[507]  & ~\main_1/preS<17>0.1 )) | ((\[617]  & (~\[541]  & \main_1/preS<17>0.1 )) | ((\[584]  & (\[582]  & \main_1/preS<12>0.1 )) | ((\[547]  & (\[507]  & \main_1/preS<17>0.1 )) | ((~\[541]  & (\[524]  & \main_1/preS<15>0.1 )) | ((\[617]  & \[555] ) | \[693] ))))))))),
  \[5]  = (\[493]  & \inreg<43> ) | (\[492]  & \inreg<51> ),
  \[584]  = ~\main_1/preS<16>0.1  & ~\main_1/preS<14>0.1 ,
  \[6]  = (\[493]  & \inreg<42> ) | (\[492]  & \inreg<50> ),
  \outreg_new<20>  = \[100] ,
  \[585]  = (~\main_1/S4_1/$S4<1>301.1  & \data<24> ) | (\main_1/S4_1/$S4<1>301.1  & ~\data<24> ),
  \[7]  = (\[493]  & \inreg<41> ) | (\[492]  & \inreg<49> ),
  \outreg_new<29>  = \[91] ,
  \[586]  = (~\main_1/S0_1/$S0<2>1.1  & \data<16> ) | (\main_1/S0_1/$S0<2>1.1  & ~\data<16> ),
  \[8]  = (\[493]  & \inreg<40> ) | (\[492]  & \inreg<48> ),
  \[587]  = (~\main_1/S0_1/$S0<3>1.1  & \data<8> ) | (\main_1/S0_1/$S0<3>1.1  & ~\data<8> ),
  \[9]  = (\[493]  & \inreg<39> ) | (\[492]  & \inreg<47> ),
  \[588]  = (~\main_1/S3_1/$S3<0>226.1  & \data<0> ) | (\main_1/S3_1/$S3<0>226.1  & ~\data<0> ),
  \[589]  = (~\main_1/S3_1/$S3<3>226.1  & \data<25> ) | (\main_1/S3_1/$S3<3>226.1  & ~\data<25> ),
  \main_1/preS<24>0.1  = (~\data<47>  & \D<12> ) | (\data<47>  & ~\D<12> ),
  \outreg_new<25>  = \[95] ,
  \outreg_new<26>  = \[94] ,
  \main_1/S0_1/$S0<2>1.1  = (~\[714]  & (\[557]  & (\main_1/preS<2>0.1  & ~\main_1/preS<1>0.1 ))) | ((\[567]  & (\[520]  & ~\main_1/preS<0>0.1 )) | ((\[566]  & (\[561]  & ~\main_1/preS<4>0.1 )) | ((~\[557]  & (\[548]  & ~\[528] )) | ((\[554]  & (~\main_1/preS<3>0.1  & ~\main_1/S0_1/$S0<1>1.1 )) | ((\[548]  & (\[537]  & \main_1/preS<2>0.1 )) | ((\[537]  & (\[536]  & \main_1/preS<1>0.1 )) | ((\[536]  & (~\main_1/preS<4>0.1  & ~\main_1/preS<3>0.1 )) | ((~\[528]  & (~\main_1/preS<4>0.1  & \main_1/preS<3>0.1 )) | ((\[714]  & \[520] ) | ((\[709]  & ~\main_1/preS<0>0.1 ) | ((\[677]  & ~\main_1/S0_1/$S0<1>1.1 ) | ((\[661]  & \main_1/preS<0>0.1 ) | \$$COND34<0>1.1 )))))))))))),
  \outreg_new<27>  = \[93] ,
  \main_1/S3_1/$S3<3>226.1  = (~\[664]  & (\[651]  & (~\[618]  & (\main_1/preS<21>0.1  & ~\$$COND233<0>226.1 )))) | ((\[669]  & (~\[628]  & (~\[535]  & \main_1/preS<19>0.1 ))) | ((\[628]  & (~\[572]  & (~\main_1/preS<19>0.1  & ~\$$COND233<0>226.1 ))) | ((\[729]  & (\[627]  & \[535] )) | ((\[729]  & (\[551]  & \[533] )) | ((\[664]  & (~\[651]  & ~\[552] )) | ((~\[628]  & (\[572]  & ~\main_1/preS<19>0.1 )) | ((\[627]  & (\[552]  & ~\[510] )) | ((\[529]  & (\main_1/preS<21>0.1  & \main_1/preS<19>0.1 )) | ((\[650]  & \[618] ) | (\$$COND238<0>226.1  | \$$COND196<0>226.1 )))))))))),
  \outreg_new<28>  = \[92] ,
  \main_1/S4_1/$S4<2>301.1  = (~\[581]  & (~\[565]  & (~\[553]  & (~\[527]  & ~\[521] )))) | ((~\[630]  & (~\[576]  & (\[553]  & ~\[527] ))) | ((\[581]  & (~\[565]  & (~\[553]  & \[526] ))) | ((\[630]  & (\[575]  & \[565] )) | ((\[630]  & (\[526]  & ~\main_1/preS<29>0.1 )) | ((\[576]  & (\[575]  & \[546] )) | ((\[565]  & (\[521]  & ~\[506] )) | ((\[565]  & (\[506]  & ~\main_1/preS<26>0.1 )) | ((\[553]  & (\[506]  & \[504] )) | ((\[546]  & (\[521]  & \main_1/preS<28>0.1 )) | ((\[540]  & (\[506]  & ~\[504] )) | (\[526]  & (~\[504]  & \main_1/preS<29>0.1 )))))))))))),
  \outreg_new<31>  = \[89] ,
  \main_1/S1_1/$S1<3>76.1  = (~\[732]  & (~\[657]  & (~\[640]  & (~\[570]  & (\[508]  & ~\main_1/preS<11>0.1 ))))) | ((~\[717]  & (\[523]  & (\main_1/preS<9>0.1  & (~\main_1/preS<8>0.1  & (~\main_1/preS<11>0.1  & ~\$$COND99<0>76.1 ))))) | ((~\[678]  & (~\[657]  & (~\[629]  & (\[571]  & ~\[538] )))) | ((~\[678]  & (~\[538]  & (~\main_1/preS<8>0.1  & (\main_1/preS<11>0.1  & \main_1/preS<10>0.1 )))) | ((\[640]  & (\[508]  & (\main_1/preS<7>0.1  & ~\main_1/preS<11>0.1 ))) | ((\[678]  & (\[657]  & \[571] )) | ((\[678]  & (~\main_1/preS<8>0.1  & ~\main_1/preS<10>0.1 )) | ((\[571]  & (\[538]  & ~\main_1/preS<6>0.1 )) | ((\[570]  & (~\main_1/preS<7>0.1  & \main_1/preS<11>0.1 )) | ((\[732]  & ~\[508] ) | ((\[724]  & \[629] ) | \$$COND70<0>76.1 )))))))))),
  \outreg_new<32>  = \[88] ,
  \$$COND34<0>1.1  = \[554]  & (\[536]  & ~\[518] ),
  \outreg_new<33>  = \[87] ,
  \[590]  = (~\main_1/S1_1/$S1<0>76.1  & \data<17> ) | (\main_1/S1_1/$S1<0>76.1  & ~\data<17> ),
  \main_1/preS<36>0.1  = (~\data<55>  & \D<15> ) | (\data<55>  & ~\D<15> ),
  \outreg_new<34>  = \[86] ,
  \[591]  = (~\main_1/S3_1/$S3<1>226.1  & \data<9> ) | (\main_1/S3_1/$S3<1>226.1  & ~\data<9> ),
  \[592]  = (~\main_1/S1_1/$S1<1>76.1  & \data<1> ) | (\main_1/S1_1/$S1<1>76.1  & ~\data<1> ),
  \[593]  = (~\main_1/S7_1/$S7<2>526.1  & \data<26> ) | (\main_1/S7_1/$S7<2>526.1  & ~\data<26> ),
  \[594]  = (~\main_1/S5_1/$S5<0>376.1  & \data<18> ) | (\main_1/S5_1/$S5<0>376.1  & ~\data<18> ),
  \outreg_new<30>  = \[90] ,
  \[595]  = (~\main_1/S5_1/$S5<1>376.1  & \data<10> ) | (\main_1/S5_1/$S5<1>376.1  & ~\data<10> ),
  \outreg_new<39>  = \[81] ,
  \[596]  = (~\main_1/S4_1/$S4<0>301.1  & \data<2> ) | (\main_1/S4_1/$S4<0>301.1  & ~\data<2> ),
  \[597]  = (~\main_1/S1_1/$S1<2>76.1  & \data<27> ) | (\main_1/S1_1/$S1<2>76.1  & ~\data<27> ),
  \[598]  = (~\main_1/S3_1/$S3<2>226.1  & \data<19> ) | (\main_1/S3_1/$S3<2>226.1  & ~\data<19> ),
  \$$COND238<0>226.1  = \[704]  & \[641] ,
  \[599]  = (~\main_1/S6_1/$S6<2>451.1  & \data<11> ) | (\main_1/S6_1/$S6<2>451.1  & ~\data<11> ),
  \outreg_new<35>  = \[85] ,
  \outreg_new<36>  = \[84] ,
  \outreg_new<37>  = \[83] ,
  \$$COND95<0>76.1  = 0,
  \outreg_new<38>  = \[82] ,
  \outreg_new<41>  = \[79] ,
  \outreg_new<42>  = \[78] ,
  \main_1/preS<20>0.1  = (~\data<45>  & \C<26> ) | (\data<45>  & ~\C<26> ),
  \outreg_new<43>  = \[77] ,
  \$$COND99<0>76.1  = \[674]  & \[570] ,
  \outreg_new<44>  = \[76] ,
  \main_1/preS<2>0.1  = (~\data<33>  & \C<10> ) | (\data<33>  & ~\C<10> ),
  \outreg_new<40>  = \[80] ,
  \outreg_new<49>  = \[71] ,
  \main_1/preS<32>0.1  = (~\data<53>  & \D<22> ) | (\data<53>  & ~\D<22> ),
  \$$COND196<0>226.1  = \[653]  & \[637] ,
  \outreg_new<45>  = \[75] ,
  \outreg_new<46>  = \[74] ,
  \outreg_new<47>  = \[73] ,
  \outreg_new<48>  = \[72] ,
  \main_1/S5_1/$S5<0>376.1  = (~\[701]  & (~\[578]  & (~\[532]  & (~\[516]  & ~\main_1/preS<31>0.1 )))) | ((~\[671]  & (~\[642]  & (~\[569]  & (~\[525]  & \main_1/preS<31>0.1 )))) | ((\[670]  & (\[525]  & ~\main_1/preS<35>0.1 )) | ((\[702]  & ~\main_1/preS<34>0.1 ) | ((\[701]  & \[516] ) | ((\[673]  & \main_1/preS<30>0.1 ) | ((\[671]  & \[635] ) | ((\[659]  & \[635] ) | ((\[625]  & ~\[532] ) | ((\[569]  & \[525] ) | ((\[532]  & ~\[505] ) | \$$COND359<0>376.1 )))))))))),
  \main_1/preS<45>0.1  = (~\data<62>  & \D<7> ) | (\data<62>  & ~\D<7> ),
  \$$COND76<0>76.1  = \[666]  & ~\[508] ,
  \$$COND484<0>526.1  = \[649]  & (\main_1/preS<47>0.1  & \main_1/preS<44>0.1 ),
  \$$COND70<0>76.1  = \[732]  & (\[622]  & ~\main_1/preS<6>0.1 ),
  \main_1/preS<18>0.1  = (~\data<43>  & \C<15> ) | (\data<43>  & ~\C<15> ),
  \main_1/preS<41>0.1  = (~\data<60>  & \D<24> ) | (\data<60>  & ~\D<24> ),
  \main_1/S4_1/$S4<1>301.1  = (\[581]  & (~\[575]  & (~\[556]  & (~\[546]  & ~\[540] )))) | ((\[576]  & (\main_1/preS<27>0.1  & ~\main_1/preS<24>0.1 )) | ((\[575]  & (\[553]  & \[521] )) | ((\[575]  & (~\main_1/preS<27>0.1  & \main_1/preS<25>0.1 )) | ((\[546]  & (~\[527]  & ~\[504] )) | ((\[546]  & (\[504]  & ~\main_1/preS<28>0.1 )) | ((~\[527]  & (\[504]  & ~\main_1/preS<29>0.1 )) | ((\[527]  & (\[521]  & ~\main_1/preS<29>0.1 )) | ((\[728]  & \[540] ) | ((\[725]  & ~\main_1/preS<25>0.1 ) | (\[703]  & \[630] )))))))))),
  \$$COND43<0>1.1  = 0,
  \main_1/S6_1/$S6<0>451.1  = (~\[713]  & (\[573]  & (\[514]  & (\main_1/preS<41>0.1  & \main_1/preS<36>0.1 )))) | ((\[667]  & (~\[522]  & (~\[514]  & \main_1/preS<41>0.1 ))) | ((\[645]  & (\[574]  & (\[573]  & \main_1/preS<39>0.1 ))) | ((~\[644]  & (~\[573]  & (\[512]  & ~\main_1/preS<40>0.1 ))) | ((~\[638]  & (\[624]  & (~\[574]  & ~\main_1/preS<39>0.1 ))) | ((~\[638]  & (~\[522]  & (~\main_1/preS<41>0.1  & \main_1/preS<36>0.1 ))) | ((\[727]  & (\[514]  & \main_1/preS<41>0.1 )) | ((\[719]  & (\[522]  & ~\main_1/preS<36>0.1 )) | ((\[667]  & (\[638]  & \main_1/preS<38>0.1 )) | ((~\[645]  & (\[631]  & ~\main_1/preS<39>0.1 )) | ((\[645]  & (\[644]  & ~\$$COND414<0>451.1 )) | ((\[573]  & (\[542]  & \[512] )) | ((\[633]  & \[631] ) | \[682] )))))))))))),
  \$$COND82<0>76.1  = 0,
  \$$COND157<0>151.1  = 0,
  \$$COND307<0>301.1  = 0,
  \[200]  = (\[503]  & \C<15> ) | ((\[502]  & \C<17> ) | ((\[501]  & \C<18> ) | ((\[500]  & \C<14> ) | ((\[499]  & \C<16> ) | ((\[498]  & \inreg<42> ) | (\[497]  & \inreg<50> )))))),
  \[201]  = (\[503]  & \C<14> ) | ((\[502]  & \C<16> ) | ((\[501]  & \C<17> ) | ((\[500]  & \C<13> ) | ((\[499]  & \C<15> ) | ((\[498]  & \inreg<50> ) | (\[497]  & \data_in<1> )))))),
  \[202]  = (\[503]  & \C<13> ) | ((\[502]  & \C<15> ) | ((\[501]  & \C<16> ) | ((\[500]  & \C<12> ) | ((\[499]  & \C<14> ) | ((\[498]  & \data_in<1> ) | (\[497]  & \inreg<1> )))))),
  \main_1/preS<14>0.1  = (~\data<41>  & \C<11> ) | (\data<41>  & ~\C<11> ),
  \[203]  = (\[503]  & \C<12> ) | ((\[502]  & \C<14> ) | ((\[501]  & \C<15> ) | ((\[500]  & \C<11> ) | ((\[499]  & \C<13> ) | ((\[498]  & \inreg<1> ) | (\[497]  & \inreg<9> )))))),
  \[204]  = (\[503]  & \C<11> ) | ((\[502]  & \C<13> ) | ((\[501]  & \C<14> ) | ((\[500]  & \C<10> ) | ((\[499]  & \C<12> ) | ((\[498]  & \inreg<9> ) | (\[497]  & \inreg<17> )))))),
  \[205]  = (\[503]  & \C<10> ) | ((\[502]  & \C<12> ) | ((\[501]  & \C<13> ) | ((\[500]  & \C<9> ) | ((\[499]  & \C<11> ) | ((\[498]  & \inreg<17> ) | (\[497]  & \inreg<25> )))))),
  \[206]  = (\[503]  & \C<9> ) | ((\[502]  & \C<11> ) | ((\[501]  & \C<12> ) | ((\[500]  & \C<8> ) | ((\[499]  & \C<10> ) | ((\[498]  & \inreg<25> ) | (\[497]  & \inreg<33> )))))),
  \main_1/preS<6>0.1  = (~\data<35>  & \C<2> ) | (\data<35>  & ~\C<2> ),
  \[207]  = (\[503]  & \C<8> ) | ((\[502]  & \C<10> ) | ((\[501]  & \C<11> ) | ((\[500]  & \C<7> ) | ((\[499]  & \C<9> ) | ((\[498]  & \inreg<33> ) | (\[497]  & \inreg<41> )))))),
  \[208]  = (\[503]  & \C<7> ) | ((\[502]  & \C<9> ) | ((\[501]  & \C<10> ) | ((\[500]  & \C<6> ) | ((\[499]  & \C<8> ) | ((\[498]  & \inreg<41> ) | (\[497]  & \inreg<49> )))))),
  \[209]  = (\[503]  & \C<6> ) | ((\[502]  & \C<8> ) | ((\[501]  & \C<9> ) | ((\[500]  & \C<5> ) | ((\[499]  & \C<7> ) | ((\[498]  & \inreg<49> ) | (\[497]  & \data_in<0> )))))),
  \$$COND65<0>76.1  = 0,
  \[210]  = (\[503]  & \C<5> ) | ((\[502]  & \C<7> ) | ((\[501]  & \C<8> ) | ((\[500]  & \C<4> ) | ((\[499]  & \C<6> ) | ((\[498]  & \data_in<0> ) | (\[497]  & \inreg<0> )))))),
  \[211]  = (\[503]  & \C<4> ) | ((\[502]  & \C<6> ) | ((\[501]  & \C<7> ) | ((\[500]  & \C<3> ) | ((\[499]  & \C<5> ) | ((\[498]  & \inreg<0> ) | (\[497]  & \inreg<8> )))))),
  \[212]  = (\[503]  & \C<3> ) | ((\[502]  & \C<5> ) | ((\[501]  & \C<6> ) | ((\[500]  & \C<2> ) | ((\[499]  & \C<4> ) | ((\[498]  & \inreg<8> ) | (\[497]  & \inreg<16> )))))),
  \[213]  = (\[503]  & \C<2> ) | ((\[502]  & \C<4> ) | ((\[501]  & \C<5> ) | ((\[500]  & \C<1> ) | ((\[499]  & \C<3> ) | ((\[498]  & \inreg<16> ) | (\[497]  & \inreg<24> )))))),
  \[214]  = (\[503]  & \C<1> ) | ((\[502]  & \C<3> ) | ((\[501]  & \C<4> ) | ((\[500]  & \C<0> ) | ((\[499]  & \C<2> ) | ((\[498]  & \inreg<24> ) | (\[497]  & \inreg<32> )))))),
  \main_1/preS<27>0.1  = (~\data<50>  & \D<8> ) | (\data<50>  & ~\D<8> ),
  \[215]  = (\[503]  & \C<0> ) | ((\[502]  & \C<2> ) | ((\[501]  & \C<3> ) | ((\[500]  & \C<27> ) | ((\[499]  & \C<1> ) | ((\[498]  & \inreg<32> ) | (\[497]  & \inreg<40> )))))),
  \C_new<23>  = \[193] ,
  \[216]  = (\[503]  & \C<27> ) | ((\[502]  & \C<1> ) | ((\[501]  & \C<2> ) | ((\[500]  & \C<26> ) | ((\[499]  & \C<0> ) | ((\[498]  & \inreg<40> ) | (\[497]  & \inreg<48> )))))),
  \C_new<24>  = \[192] ,
  \$$COND281<0>301.1  = 0,
  \[217]  = (\[503]  & \D<26> ) | ((\[502]  & \D<0> ) | ((\[501]  & \D<1> ) | ((\[500]  & \D<25> ) | ((\[499]  & \D<27> ) | ((\[498]  & \inreg<54> ) | (\[497]  & \data_in<3> )))))),
  \C_new<21>  = \[195] ,
  \main_1/S0_1/$S0<3>1.1  = (~\[714]  & (\[562]  & (\[554]  & (~\[536]  & ~\main_1/preS<1>0.1 )))) | ((~\[566]  & (~\[548]  & (\[537]  & \[528] ))) | ((~\[562]  & (~\[554]  & (~\[520]  & ~\main_1/preS<1>0.1 ))) | ((~\[554]  & (~\[528]  & (~\[520]  & \main_1/preS<1>0.1 ))) | ((\[706]  & (~\[562]  & \[554] )) | ((\[567]  & (~\[557]  & \[536] )) | ((\[567]  & (\[557]  & \main_1/preS<2>0.1 )) | ((\[562]  & (\[548]  & \[520] )) | ((\[557]  & (\[536]  & ~\main_1/preS<1>0.1 )) | ((\[554]  & (\[536]  & \main_1/preS<3>0.1 )) | \[661] ))))))))),
  \[218]  = (\[503]  & \D<25> ) | ((\[502]  & \D<27> ) | ((\[501]  & \D<0> ) | ((\[500]  & \D<24> ) | ((\[499]  & \D<26> ) | ((\[498]  & \data_in<3> ) | (\[497]  & \inreg<3> )))))),
  \C_new<22>  = \[194] ,
  \main_1/preS<10>0.1  = (~\data<39>  & \C<20> ) | (\data<39>  & ~\C<20> ),
  \[219]  = (\[503]  & \D<24> ) | ((\[502]  & \D<26> ) | ((\[501]  & \D<27> ) | ((\[500]  & \D<23> ) | ((\[499]  & \D<25> ) | ((\[498]  & \inreg<3> ) | (\[497]  & \inreg<11> )))))),
  \$$COND311<0>301.1  = \[581]  & ~\[527] ,
  \C_new<20>  = \[196] ,
  \main_1/preS<39>0.1  = (~\data<58>  & \D<27> ) | (\data<58>  & ~\D<27> ),
  \data_new<4>  = \[180] ,
  \[220]  = (\[503]  & \D<23> ) | ((\[502]  & \D<25> ) | ((\[501]  & \D<26> ) | ((\[500]  & \D<22> ) | ((\[499]  & \D<24> ) | ((\[498]  & \inreg<11> ) | (\[497]  & \inreg<19> )))))),
  \data_new<3>  = \[181] ,
  \[600]  = (~\main_1/S5_1/$S5<3>376.1  & \data<3> ) | (\main_1/S5_1/$S5<3>376.1  & ~\data<3> ),
  \[221]  = (\[503]  & \D<22> ) | ((\[502]  & \D<24> ) | ((\[501]  & \D<25> ) | ((\[500]  & \D<21> ) | ((\[499]  & \D<23> ) | ((\[498]  & \inreg<19> ) | (\[497]  & \data_in<4> )))))),
  \C_new<27>  = \[189] ,
  \data_new<2>  = \[182] ,
  \[601]  = (~\main_1/S5_1/$S5<2>376.1  & \data<28> ) | (\main_1/S5_1/$S5<2>376.1  & ~\data<28> ),
  \[222]  = (\[503]  & \D<21> ) | ((\[502]  & \D<23> ) | ((\[501]  & \D<24> ) | ((\[500]  & \D<20> ) | ((\[499]  & \D<22> ) | ((\[498]  & \data_in<4> ) | (\[497]  & \inreg<4> )))))),
  \data_new<1>  = \[183] ,
  \[602]  = (~\main_1/S7_1/$S7<0>526.1  & \data<20> ) | (\main_1/S7_1/$S7<0>526.1  & ~\data<20> ),
  \[223]  = (\[503]  & \D<20> ) | ((\[502]  & \D<22> ) | ((\[501]  & \D<23> ) | ((\[500]  & \D<19> ) | ((\[499]  & \D<21> ) | ((\[498]  & \inreg<4> ) | (\[497]  & \inreg<12> )))))),
  \C_new<25>  = \[191] ,
  \data_new<0>  = \[184] ,
  \[603]  = (~\main_1/S1_1/$S1<3>76.1  & \data<12> ) | (\main_1/S1_1/$S1<3>76.1  & ~\data<12> ),
  \[224]  = (\[503]  & \D<19> ) | ((\[502]  & \D<21> ) | ((\[501]  & \D<22> ) | ((\[500]  & \D<18> ) | ((\[499]  & \D<20> ) | ((\[498]  & \inreg<12> ) | (\[497]  & \inreg<20> )))))),
  \C_new<26>  = \[190] ,
  \[604]  = (~\main_1/S7_1/$S7<3>526.1  & \data<4> ) | (\main_1/S7_1/$S7<3>526.1  & ~\data<4> ),
  \[225]  = (\[503]  & \D<18> ) | ((\[502]  & \D<20> ) | ((\[501]  & \D<21> ) | ((\[500]  & \D<17> ) | ((\[499]  & \D<19> ) | ((\[498]  & \inreg<20> ) | (\[497]  & \inreg<28> )))))),
  \C_new<13>  = \[203] ,
  \[605]  = (~\main_1/S2_1/$S2<1>151.1  & \data<29> ) | (\main_1/S2_1/$S2<1>151.1  & ~\data<29> ),
  \[226]  = (\[503]  & \D<17> ) | ((\[502]  & \D<19> ) | ((\[501]  & \D<20> ) | ((\[500]  & \D<16> ) | ((\[499]  & \D<18> ) | ((\[498]  & \inreg<28> ) | (\[497]  & \inreg<36> )))))),
  \C_new<14>  = \[202] ,
  \[606]  = (~\main_1/S6_1/$S6<1>451.1  & \data<21> ) | (\main_1/S6_1/$S6<1>451.1  & ~\data<21> ),
  \[227]  = (\[503]  & \D<16> ) | ((\[502]  & \D<18> ) | ((\[501]  & \D<19> ) | ((\[500]  & \D<15> ) | ((\[499]  & \D<17> ) | ((\[498]  & \inreg<36> ) | (\[497]  & \inreg<44> )))))),
  \C_new<11>  = \[205] ,
  \[607]  = (~\main_1/S4_1/$S4<2>301.1  & \data<13> ) | (\main_1/S4_1/$S4<2>301.1  & ~\data<13> ),
  \[228]  = (\[503]  & \D<15> ) | ((\[502]  & \D<17> ) | ((\[501]  & \D<18> ) | ((\[500]  & \D<14> ) | ((\[499]  & \D<16> ) | ((\[498]  & \inreg<44> ) | (\[497]  & \inreg<52> )))))),
  \C_new<12>  = \[204] ,
  \[608]  = (~\main_1/S2_1/$S2<0>151.1  & \data<5> ) | (\main_1/S2_1/$S2<0>151.1  & ~\data<5> ),
  \$$COND371<0>376.1  = \[659]  & \[643] ,
  \[229]  = (\[503]  & \D<14> ) | ((\[502]  & \D<16> ) | ((\[501]  & \D<17> ) | ((\[500]  & \D<13> ) | ((\[499]  & \D<15> ) | ((\[498]  & \inreg<52> ) | (\[497]  & \data_in<5> )))))),
  \[609]  = (~\main_1/S0_1/$S0<0>1.1  & \data<30> ) | (\main_1/S0_1/$S0<0>1.1  & ~\data<30> ),
  \C_new<10>  = \[206] ,
  \data_new<9>  = \[175] ,
  \main_1/S2_1/$S2<3>151.1  = (~\[676]  & (~\[663]  & (~\[617]  & (~\[558]  & ~\[524] )))) | ((~\[663]  & (~\[530]  & (\[519]  & (\main_1/preS<15>0.1  & ~\main_1/S2_1/$S2<1>151.1 )))) | ((~\[676]  & (~\[519]  & (\main_1/preS<16>0.1  & \main_1/preS<15>0.1 ))) | ((~\[507]  & (~\main_1/preS<16>0.1  & (~\main_1/preS<15>0.1  & ~\main_1/preS<12>0.1 ))) | ((\[676]  & (~\[519]  & \main_1/S2_1/$S2<1>151.1 )) | ((\[672]  & (\[507]  & ~\main_1/preS<12>0.1 )) | ((\[656]  & (\[555]  & \main_1/S2_1/$S2<1>151.1 )) | ((\[623]  & (\[530]  & \[507] )) | ((\[582]  & (~\[541]  & \[530] )) | ((\[558]  & (\main_1/preS<12>0.1  & \main_1/S2_1/$S2<1>151.1 )) | (\[617]  & \[530] )))))))))),
  \main_1/preS<23>0.1  = (~\data<48>  & \C<1> ) | (\data<48>  & ~\C<1> ),
  \data_new<8>  = \[176] ,
  \data_new<7>  = \[177] ,
  \main_1/S5_1/$S5<2>376.1  = (~\[670]  & (~\[632]  & (~\[578]  & (~\[532]  & (\[505]  & ~\main_1/S5_1/$S5<3>376.1 ))))) | ((~\[643]  & (~\[642]  & (~\[620]  & (~\main_1/preS<32>0.1  & \main_1/S5_1/$S5<3>376.1 )))) | ((\[659]  & (~\[578]  & (\[569]  & ~\[532] ))) | ((\[642]  & (~\[505]  & (~\main_1/preS<35>0.1  & \main_1/S5_1/$S5<3>376.1 ))) | ((~\[505]  & (\main_1/preS<35>0.1  & (~\main_1/preS<34>0.1  & ~\main_1/S5_1/$S5<3>376.1 ))) | ((\[702]  & (\[632]  & \[578] )) | ((\[670]  & (~\[620]  & ~\main_1/preS<35>0.1 )) | ((~\[659]  & (\[643]  & \[505] )) | ((\[659]  & (~\[569]  & \main_1/preS<34>0.1 )) | ((\[702]  & \[673] ) | (\[620]  & ~\[505] )))))))))),
  \data_new<6>  = \[178] ,
  \data_new<5>  = \[179] ,
  \C_new<19>  = \[197] ,
  \[230]  = (\[503]  & \D<13> ) | ((\[502]  & \D<15> ) | ((\[501]  & \D<16> ) | ((\[500]  & \D<12> ) | ((\[499]  & \D<14> ) | ((\[498]  & \data_in<5> ) | (\[497]  & \inreg<5> )))))),
  \[610]  = (~\main_1/S0_1/$S0<1>1.1  & \data<22> ) | (\main_1/S0_1/$S0<1>1.1  & ~\data<22> ),
  \[231]  = (\[503]  & \D<12> ) | ((\[502]  & \D<14> ) | ((\[501]  & \D<15> ) | ((\[500]  & \D<11> ) | ((\[499]  & \D<13> ) | ((\[498]  & \inreg<5> ) | (\[497]  & \inreg<13> )))))),
  \C_new<17>  = \[199] ,
  \[611]  = (~\main_1/S7_1/$S7<1>526.1  & \data<14> ) | (\main_1/S7_1/$S7<1>526.1  & ~\data<14> ),
  \[232]  = (\[503]  & \D<11> ) | ((\[502]  & \D<13> ) | ((\[501]  & \D<14> ) | ((\[500]  & \D<10> ) | ((\[499]  & \D<12> ) | ((\[498]  & \inreg<13> ) | (\[497]  & \inreg<21> )))))),
  \C_new<18>  = \[198] ,
  \main_1/preS<35>0.1  = (~\data<56>  & \D<19> ) | (\data<56>  & ~\D<19> ),
  \[612]  = (~\main_1/S6_1/$S6<0>451.1  & \data<6> ) | (\main_1/S6_1/$S6<0>451.1  & ~\data<6> ),
  \[233]  = (\[503]  & \D<10> ) | ((\[502]  & \D<12> ) | ((\[501]  & \D<13> ) | ((\[500]  & \D<9> ) | ((\[499]  & \D<11> ) | ((\[498]  & \inreg<21> ) | (\[497]  & \inreg<29> )))))),
  \C_new<15>  = \[201] ,
  \[613]  = (~\main_1/S6_1/$S6<3>451.1  & \data<31> ) | (\main_1/S6_1/$S6<3>451.1  & ~\data<31> ),
  \[234]  = (\[503]  & \D<9> ) | ((\[502]  & \D<11> ) | ((\[501]  & \D<12> ) | ((\[500]  & \D<8> ) | ((\[499]  & \D<10> ) | ((\[498]  & \inreg<29> ) | (\[497]  & \inreg<37> )))))),
  \C_new<16>  = \[200] ,
  \[614]  = (~\main_1/S2_1/$S2<3>151.1  & \data<23> ) | (\main_1/S2_1/$S2<3>151.1  & ~\data<23> ),
  \[235]  = (\[503]  & \D<8> ) | ((\[502]  & \D<10> ) | ((\[501]  & \D<11> ) | ((\[500]  & \D<7> ) | ((\[499]  & \D<9> ) | ((\[498]  & \inreg<37> ) | (\[497]  & \inreg<45> )))))),
  \D_new<13>  = \[231] ,
  \[615]  = (~\main_1/S2_1/$S2<2>151.1  & \data<15> ) | (\main_1/S2_1/$S2<2>151.1  & ~\data<15> ),
  \[236]  = (\[503]  & \D<7> ) | ((\[502]  & \D<9> ) | ((\[501]  & \D<10> ) | ((\[500]  & \D<6> ) | ((\[499]  & \D<8> ) | ((\[498]  & \inreg<45> ) | (\[497]  & \inreg<53> )))))),
  \D_new<14>  = \[230] ,
  \[616]  = (~\main_1/S4_1/$S4<3>301.1  & \data<7> ) | (\main_1/S4_1/$S4<3>301.1  & ~\data<7> ),
  \[237]  = (\[503]  & \D<6> ) | ((\[502]  & \D<8> ) | ((\[501]  & \D<9> ) | ((\[500]  & \D<5> ) | ((\[499]  & \D<7> ) | ((\[498]  & \inreg<53> ) | (\[497]  & \data_in<6> )))))),
  \D_new<11>  = \[233] ,
  \[617]  = (\[547]  & ~\main_1/preS<14>0.1 ) | (~\[509]  & ~\main_1/preS<16>0.1 ),
  \[238]  = (\[503]  & \D<5> ) | ((\[502]  & \D<7> ) | ((\[501]  & \D<8> ) | ((\[500]  & \D<4> ) | ((\[499]  & \D<6> ) | ((\[498]  & \data_in<6> ) | (\[497]  & \inreg<6> )))))),
  \D_new<12>  = \[232] ,
  \[618]  = ~\main_1/preS<20>0.1  & \main_1/preS<18>0.1 ,
  \[239]  = (\[503]  & \D<4> ) | ((\[502]  & \D<6> ) | ((\[501]  & \D<7> ) | ((\[500]  & \D<3> ) | ((\[499]  & \D<5> ) | ((\[498]  & \inreg<6> ) | (\[497]  & \inreg<14> )))))),
  \[619]  = \main_1/preS<35>0.1  & \main_1/preS<31>0.1 ,
  \D_new<10>  = \[234] ,
  \data_new<63>  = \[121] ,
  \data_new<61>  = \[123] ,
  \data_new<62>  = \[122] ,
  \D_new<19>  = \[225] ,
  \data_new<60>  = \[124] ,
  \[240]  = (\[503]  & \D<3> ) | ((\[502]  & \D<5> ) | ((\[501]  & \D<6> ) | ((\[500]  & \D<2> ) | ((\[499]  & \D<4> ) | ((\[498]  & \inreg<14> ) | (\[497]  & \inreg<22> )))))),
  \[620]  = \[525]  & ~\main_1/preS<35>0.1 ,
  \[241]  = (\[503]  & \D<2> ) | ((\[502]  & \D<4> ) | ((\[501]  & \D<5> ) | ((\[500]  & \D<1> ) | ((\[499]  & \D<3> ) | ((\[498]  & \inreg<22> ) | (\[497]  & \inreg<30> )))))),
  \D_new<17>  = \[227] ,
  \[621]  = \[534]  & ~\main_1/preS<46>0.1 ,
  \[242]  = (\[503]  & \D<1> ) | ((\[502]  & \D<3> ) | ((\[501]  & \D<4> ) | ((\[500]  & \D<0> ) | ((\[499]  & \D<2> ) | ((\[498]  & \inreg<30> ) | (\[497]  & \inreg<38> )))))),
  \D_new<18>  = \[226] ,
  \[622]  = ~\main_1/preS<9>0.1  & ~\main_1/preS<7>0.1 ,
  \[243]  = (\[503]  & \D<0> ) | ((\[502]  & \D<2> ) | ((\[501]  & \D<3> ) | ((\[500]  & \D<27> ) | ((\[499]  & \D<1> ) | ((\[498]  & \inreg<38> ) | (\[497]  & \inreg<46> )))))),
  \D_new<15>  = \[229] ,
  \[623]  = ~\[509]  & \main_1/preS<16>0.1 ,
  \[244]  = (\[503]  & \D<27> ) | ((\[502]  & \D<1> ) | ((\[501]  & \D<2> ) | ((\[500]  & \D<26> ) | ((\[499]  & \D<0> ) | ((\[498]  & \inreg<46> ) | (\[497]  & \inreg<54> )))))),
  \D_new<16>  = \[228] ,
  \[624]  = \main_1/preS<38>0.1  & ~\main_1/preS<36>0.1 ,
  \[245]  = (~\generate_key_1/freeze<0>605.1  & \encrypt_mode<0> ) | (\generate_key_1/freeze<0>605.1  & \encrypt<0> ),
  \D_new<23>  = \[221] ,
  \[625]  = \[569]  & ~\main_1/preS<32>0.1 ,
  \main_1/preS<1>0.1  = (~\data<32>  & \C<16> ) | (\data<32>  & ~\C<16> ),
  \D_new<24>  = \[220] ,
  \[626]  = \main_1/preS<19>0.1  & ~\main_1/preS<18>0.1 ,
  \D_new<21>  = \[223] ,
  \[627]  = \main_1/preS<23>0.1  & ~\main_1/preS<22>0.1 ,
  \D_new<22>  = \[222] ,
  \[628]  = \main_1/preS<20>0.1  & \main_1/preS<18>0.1 ,
  \main_1/preS<31>0.1  = (~\data<52>  & \D<11> ) | (\data<52>  & ~\D<11> ),
  \[629]  = \main_1/preS<6>0.1  & ~\main_1/preS<10>0.1 ,
  \D_new<20>  = \[224] ,
  \data_new<53>  = \[131] ,
  \data_new<54>  = \[130] ,
  \data_new<51>  = \[133] ,
  \data_new<52>  = \[132] ,
  \main_1/S6_1/$S6<2>451.1  = (~\[634]  & (~\[542]  & (\[514]  & (~\main_1/preS<38>0.1  & ~\main_1/preS<36>0.1 )))) | ((~\[667]  & (\[550]  & (\main_1/preS<40>0.1  & \main_1/preS<38>0.1 ))) | ((\[667]  & (\[550]  & (~\main_1/preS<40>0.1  & \main_1/preS<38>0.1 ))) | ((~\[727]  & (\[638]  & ~\main_1/preS<38>0.1 )) | ((\[645]  & (~\main_1/preS<39>0.1  & ~\main_1/preS<37>0.1 )) | ((\[631]  & (\main_1/preS<40>0.1  & \main_1/preS<36>0.1 )) | ((\[624]  & (\[542]  & \main_1/preS<37>0.1 )) | ((\[722]  & \main_1/preS<36>0.1 ) | ((\[719]  & ~\main_1/preS<37>0.1 ) | ((\[644]  & \[639] ) | (\[634]  & \main_1/preS<36>0.1 )))))))))),
  \data_new<50>  = \[134] ,
  \[630]  = \main_1/preS<26>0.1  & \main_1/preS<25>0.1 ,
  \D_new<27>  = \[217] ,
  \[631]  = \[550]  & ~\main_1/preS<38>0.1 ,
  \[632]  = \main_1/preS<32>0.1  & \main_1/preS<30>0.1 ,
  \D_new<25>  = \[219] ,
  \[633]  = \[512]  & \main_1/preS<40>0.1 ,
  \D_new<26>  = \[218] ,
  \[634]  = (\[573]  & (\main_1/preS<41>0.1  & \main_1/preS<40>0.1 )) | ((\[638]  & \main_1/preS<37>0.1 ) | (\[574]  & ~\[522] )),
  \data_new<59>  = \[125] ,
  \[635]  = \[545]  & ~\main_1/preS<33>0.1 ,
  \[636]  = \[532]  & ~\main_1/preS<35>0.1 ,
  \data_new<57>  = \[127] ,
  \[637]  = \[533]  & \main_1/preS<22>0.1 ,
  \data_new<58>  = \[126] ,
  \[638]  = ~\[514]  & ~\main_1/preS<41>0.1 ,
  \data_new<55>  = \[129] ,
  \[639]  = \[542]  & \[512] ,
  \data_new<56>  = \[128] ,
  \main_1/preS<44>0.1  = (~\data<61>  & \D<21> ) | (\data<61>  & ~\D<21> ),
  \main_1/S7_1/$S7<0>526.1  = (~\[583]  & (~\[559]  & (\[549]  & \main_1/S7_1/$S7<2>526.1 ))) | ((\[583]  & (~\main_1/preS<44>0.1  & (\main_1/preS<43>0.1  & ~\main_1/S7_1/$S7<2>526.1 ))) | ((~\[517]  & (~\main_1/preS<47>0.1  & (\main_1/preS<44>0.1  & \main_1/S7_1/$S7<2>526.1 ))) | ((~\[517]  & (\main_1/preS<44>0.1  & (~\main_1/preS<43>0.1  & ~\main_1/S7_1/$S7<2>526.1 ))) | ((\[517]  & (\main_1/preS<46>0.1  & (~\main_1/preS<44>0.1  & ~\main_1/preS<43>0.1 ))) | ((~\main_1/preS<45>0.1  & (~\main_1/preS<44>0.1  & (~\main_1/preS<43>0.1  & \main_1/S7_1/$S7<2>526.1 ))) | ((\[649]  & (~\main_1/preS<45>0.1  & ~\main_1/preS<44>0.1 )) | ((\[621]  & (~\main_1/preS<43>0.1  & ~\main_1/preS<42>0.1 )) | ((\[621]  & (\main_1/preS<43>0.1  & \main_1/preS<42>0.1 )) | ((\[559]  & (\main_1/preS<44>0.1  & \main_1/preS<43>0.1 )) | ((~\[511]  & (~\main_1/preS<47>0.1  & ~\main_1/S7_1/$S7<2>526.1 )) | ((\[711]  & \main_1/preS<47>0.1 ) | (\[662]  & \main_1/preS<47>0.1 )))))))))))),
  \[640]  = ~\[523]  & \main_1/preS<8>0.1 ,
  \main_1/S1_1/$S1<1>76.1  = (~\[710]  & (~\[640]  & (\[515]  & (~\[508]  & ~\main_1/preS<11>0.1 )))) | ((\[710]  & (~\[678]  & (~\[622]  & ~\$$COND76<0>76.1 ))) | ((\[732]  & (\main_1/preS<7>0.1  & \main_1/preS<6>0.1 )) | ((\[640]  & (\[571]  & \main_1/preS<7>0.1 )) | ((\[640]  & (\[538]  & ~\main_1/preS<11>0.1 )) | ((\[622]  & (\[544]  & ~\[515] )) | ((\[622]  & (\[515]  & ~\main_1/preS<10>0.1 )) | ((\[571]  & (~\main_1/preS<7>0.1  & \main_1/preS<10>0.1 )) | ((\[544]  & (~\[515]  & \main_1/preS<9>0.1 )) | ((\[678]  & ~\[515] ) | ((\[647]  & \[629] ) | ((\[570]  & \[538] ) | \$$COND70<0>76.1 ))))))))))),
  \[641]  = ~\main_1/preS<23>0.1  & \main_1/preS<22>0.1 ,
  \[642]  = ~\main_1/preS<34>0.1  & ~\main_1/preS<33>0.1 ,
  \[643]  = \[545]  & \main_1/preS<33>0.1 ,
  \[644]  = ~\main_1/preS<38>0.1  & \main_1/preS<37>0.1 ,
  \[645]  = ~\main_1/preS<40>0.1  & ~\main_1/preS<36>0.1 ,
  \[646]  = \[543]  & ~\main_1/preS<7>0.1 ,
  \[647]  = ~\[508]  & \main_1/preS<11>0.1 ,
  \[648]  = \count<0>  | \count<3> ,
  \$$COND225<0>226.1  = \[627]  & (\[626]  & \[551] ),
  \$$COND354<0>376.1  = \[619]  & (\[532]  & ~\[516] ),
  \$$COND244<0>226.1  = \[618]  & (\[572]  & ~\main_1/preS<19>0.1 ),
  \[649]  = ~\[517]  & \main_1/preS<43>0.1 ,
  \main_1/preS<17>0.1  = (~\data<44>  & \C<7> ) | (\data<44>  & ~\C<7> ),
  \[650]  = \[533]  & ~\main_1/preS<22>0.1 ,
  \main_1/S5_1/$S5<1>376.1  = (\[643]  & (~\main_1/preS<31>0.1  & ~\main_1/preS<30>0.1 )) | ((\[642]  & (\[619]  & \[516] )) | ((\[642]  & (\[539]  & ~\main_1/preS<30>0.1 )) | ((\[635]  & (\[632]  & ~\main_1/preS<31>0.1 )) | ((\[632]  & (\[525]  & ~\main_1/preS<31>0.1 )) | ((\[620]  & (\[505]  & \main_1/preS<31>0.1 )) | ((\[619]  & (\[578]  & ~\[516] )) | ((\[578]  & (\[539]  & \main_1/preS<30>0.1 )) | ((\[525]  & (~\[505]  & \main_1/preS<35>0.1 )) | ((\[673]  & ~\main_1/preS<32>0.1 ) | ((\[670]  & \[635] ) | ((\[643]  & ~\[505] ) | ((\[636]  & ~\[516] ) | ((\[625]  & \main_1/preS<34>0.1 ) | (\$$COND371<0>376.1  | (\$$COND354<0>376.1  | (\$$COND365<0>376.1  | (\$$COND359<0>376.1  | (\$$COND358<0>376.1  | \$$COND328<0>376.1 )))))))))))))))))),
  \main_1/preS<40>0.1  = (~\data<59>  & \D<5> ) | (\data<59>  & ~\D<5> ),
  \[651]  = ~\main_1/preS<23>0.1  & ~\main_1/preS<22>0.1 ,
  \main_1/preS<9>0.1  = (~\data<38>  & \C<5> ) | (\data<38>  & ~\C<5> ),
  \[652]  = \[534]  & ~\main_1/preS<43>0.1 ,
  \[653]  = \[535]  & ~\main_1/preS<21>0.1 ,
  \[654]  = \[535]  & \main_1/preS<21>0.1 ,
  \[655]  = ~\main_1/preS<46>0.1  & ~\main_1/preS<44>0.1 ,
  \[656]  = \main_1/preS<15>0.1  & ~\main_1/preS<13>0.1 ,
  \[657]  = ~\main_1/preS<6>0.1  & \main_1/preS<10>0.1 ,
  \main_1/S3_1/$S3<0>226.1  = (\[651]  & (\[618]  & \main_1/preS<21>0.1 )) | ((\[579]  & (~\main_1/preS<23>0.1  & ~\main_1/preS<21>0.1 )) | ((\[572]  & (\[535]  & \main_1/preS<19>0.1 )) | ((\[551]  & (\[529]  & ~\main_1/preS<18>0.1 )) | ((\[726]  & ~\main_1/preS<20>0.1 ) | ((\[669]  & \main_1/preS<19>0.1 ) | ((\[668]  & \[654] ) | ((\[664]  & \[552] ) | ((\[654]  & \[641] ) | ((\[653]  & \[533] ) | ((\[650]  & \[551] ) | ((\[637]  & \[628] ) | ((\[628]  & \[572] ) | ((\[579]  & ~\main_1/preS<22>0.1 ) | (\$$COND254<0>226.1  | (\$$COND249<0>226.1  | (\$$COND244<0>226.1  | (\$$COND216<0>226.1  | \$$COND210<0>226.1 ))))))))))))))))),
  \main_1/S4_1/$S4<3>301.1  = (~\[728]  & (~\[576]  & (\[546]  & (\[527]  & ~\[521] )))) | ((~\[660]  & (~\[630]  & (~\[581]  & (~\main_1/preS<29>0.1  & ~\main_1/S4_1/$S4<0>301.1 )))) | ((~\[703]  & (\[581]  & (\main_1/preS<29>0.1  & \main_1/preS<24>0.1 ))) | ((\[576]  & (~\main_1/preS<27>0.1  & (\main_1/preS<24>0.1  & \main_1/S4_1/$S4<0>301.1 ))) | ((\[728]  & (~\[546]  & ~\[540] )) | ((\[703]  & (~\$$COND311<0>301.1  & ~\main_1/preS<26>0.1 )) | ((\[581]  & (\[565]  & \[556] )) | ((~\[576]  & (\[540]  & ~\[527] )) | ((\[526]  & (\main_1/preS<27>0.1  & \main_1/preS<26>0.1 )) | ((\[660]  & \main_1/preS<25>0.1 ) | \[658] ))))))))),
  \[658]  = ~\[527]  & \[521] ,
  \[659]  = \[531]  & \main_1/preS<32>0.1 ,
  \[660]  = \[556]  & \[540] ,
  \[661]  = \[566]  & \[520] ,
  \$$COND520<0>0.1  = \count<3>  & (\count<2>  & (\count<1>  & \count<0> )),
  \[662]  = \[564]  & \[513] ,
  \main_1/S0_1/$S0<0>1.1  = (~\[554]  & (~\[520]  & (\main_1/preS<3>0.1  & (~\main_1/preS<0>0.1  & ~\main_1/S0_1/$S0<3>1.1 )))) | ((~\[661]  & (\[536]  & (\main_1/preS<5>0.1  & \main_1/preS<1>0.1 ))) | ((\[562]  & (~\[536]  & (\[520]  & \main_1/S0_1/$S0<3>1.1 ))) | ((\[548]  & (~\main_1/preS<4>0.1  & (\main_1/preS<0>0.1  & \main_1/S0_1/$S0<3>1.1 ))) | ((\[706]  & (\[561]  & \[537] )) | ((~\[562]  & (\[548]  & \[537] )) | ((\[554]  & (\main_1/preS<1>0.1  & \main_1/preS<0>0.1 )) | ((\[537]  & (\[536]  & ~\main_1/S0_1/$S0<3>1.1 )) | ((~\[518]  & (~\main_1/preS<4>0.1  & ~\main_1/preS<0>0.1 )) | ((\[706]  & \main_1/preS<5>0.1 ) | ((\[567]  & ~\[562] ) | (\[567]  & \[554] ))))))))))),
  \[663]  = \[547]  & ~\main_1/preS<13>0.1 ,
  \main_1/preS<13>0.1  = (~\data<40>  & \C<18> ) | (\data<40>  & ~\C<18> ),
  \[664]  = \[626]  & \main_1/preS<20>0.1 ,
  \[665]  = \[549]  & \main_1/preS<46>0.1 ,
  \[666]  = \[568]  & \[544] ,
  \[667]  = ~\main_1/preS<39>0.1  & \main_1/preS<36>0.1 ,
  \$$COND414<0>451.1  = \[645]  & (\[631]  & ~\main_1/preS<39>0.1 ),
  \main_1/preS<5>0.1  = (~\data<36>  & \C<4> ) | (\data<36>  & ~\C<4> ),
  \[668]  = \main_1/preS<23>0.1  & ~\main_1/preS<19>0.1 ,
  \[669]  = \[552]  & ~\main_1/preS<23>0.1 ,
  \[670]  = ~\[516]  & \main_1/preS<31>0.1 ,
  \[671]  = ~\main_1/preS<32>0.1  & \main_1/preS<30>0.1 ,
  \main_1/S6_1/$S6<1>451.1  = (~\main_1/preS<41>0.1  & (\main_1/preS<39>0.1  & (\main_1/preS<37>0.1  & \main_1/S6_1/$S6<2>451.1 ))) | ((\[722]  & (~\main_1/preS<39>0.1  & ~\main_1/preS<36>0.1 )) | ((\[667]  & (\[574]  & \main_1/S6_1/$S6<2>451.1 )) | ((\[644]  & (\[542]  & ~\main_1/preS<39>0.1 )) | ((\[644]  & (\[512]  & \main_1/S6_1/$S6<2>451.1 )) | ((\[624]  & (\[577]  & \main_1/preS<41>0.1 )) | ((\[550]  & (~\main_1/preS<39>0.1  & ~\main_1/preS<36>0.1 )) | ((~\[514]  & (\main_1/preS<36>0.1  & ~\main_1/S6_1/$S6<2>451.1 )) | ((\[727]  & \main_1/preS<39>0.1 ) | ((\[720]  & \main_1/preS<37>0.1 ) | ((\[716]  & \main_1/preS<38>0.1 ) | ((\[713]  & \main_1/preS<38>0.1 ) | ((\[639]  & ~\main_1/preS<37>0.1 ) | (\[682]  | \$$COND445<0>451.1 ))))))))))))),
  \[672]  = \[558]  & \main_1/preS<16>0.1 ,
  \[673]  = \[539]  & \[532] ,
  \[674]  = \[538]  & ~\main_1/preS<11>0.1 ,
  \main_1/S1_1/$S1<0>76.1  = (~\[666]  & (\[538]  & (~\main_1/preS<8>0.1  & \main_1/preS<10>0.1 ))) | ((\[629]  & (~\main_1/preS<9>0.1  & (\main_1/preS<7>0.1  & ~\main_1/preS<11>0.1 ))) | ((\[717]  & (\main_1/preS<8>0.1  & \main_1/preS<7>0.1 )) | ((\[674]  & (\main_1/preS<8>0.1  & ~\main_1/preS<10>0.1 )) | ((\[622]  & (~\main_1/preS<6>0.1  & \main_1/S1_1/$S1<3>76.1 )) | ((\[568]  & (~\main_1/preS<9>0.1  & ~\main_1/preS<11>0.1 )) | ((\[543]  & (\main_1/preS<8>0.1  & \main_1/S1_1/$S1<3>76.1 )) | ((\[674]  & \main_1/preS<6>0.1 ) | ((\[647]  & ~\main_1/S1_1/$S1<3>76.1 ) | ((\[646]  & ~\main_1/preS<10>0.1 ) | ((\[640]  & ~\[508] ) | ((\[570]  & \[543] ) | \$$COND76<0>76.1 ))))))))))),
  \[675]  = \[551]  & \main_1/preS<18>0.1 ,
  \main_1/preS<26>0.1  = (~\data<49>  & \D<2> ) | (\data<49>  & ~\D<2> ),
  \[676]  = \main_1/preS<14>0.1  & \main_1/preS<13>0.1 ,
  \[677]  = \[520]  & ~\main_1/preS<2>0.1 ,
  \[678]  = \[543]  & \main_1/preS<7>0.1 ,
  \[679]  = 0,
  \D_new<7>  = \[237] ,
  \C_new<6>  = \[210] ,
  \D_new<8>  = \[236] ,
  \C_new<5>  = \[211] ,
  \D_new<5>  = \[239] ,
  \C_new<8>  = \[208] ,
  \main_1/preS<38>0.1  = (~\data<57>  & \D<10> ) | (\data<57>  & ~\D<10> ),
  \D_new<6>  = \[238] ,
  \C_new<7>  = \[209] ,
  \C_new<9>  = \[207] ,
  \[490]  = ~\$$COND521<0>601.1  & ~\reset<0> ,
  \D_new<9>  = \[235] ,
  \[491]  = \[490]  & ~\generate_key_1/freeze<0>605.1 ,
  \[492]  = ~\count<0> ,
  \[682]  = (\[644]  & (\[638]  & \main_1/preS<36>0.1 )) | \$$COND391<0>451.1 ,
  \[493]  = ~\$$COND520<0>0.1  & \count<0> ,
  \D_new<0>  = \[244] ,
  \[494]  = \$$COND521<0>601.1  & ~\reset<0> ,
  \C_new<0>  = \[216] ,
  \[495]  = \[491]  & ~\encrypt_mode<0> ,
  \[496]  = \[491]  & \encrypt_mode<0> ,
  \D_new<3>  = \[241] ,
  \C_new<2>  = \[214] ,
  \[497]  = \[494]  & ~\encrypt<0> ,
  \D_new<4>  = \[240] ,
  \C_new<1>  = \[215] ,
  \[498]  = \[494]  & \encrypt<0> ,
  \$$COND358<0>376.1  = \[705]  & \[636] ,
  \D_new<1>  = \[243] ,
  \C_new<4>  = \[212] ,
  \[499]  = \[490]  & \generate_key_1/freeze<0>605.1 ,
  \D_new<2>  = \[242] ,
  \C_new<3>  = \[213] ,
  \main_1/preS<22>0.1  = (~\data<47>  & \C<12> ) | (\data<47>  & ~\C<12> ),
  \generate_key_1/freeze<0>605.1  = (\$$COND520<0>0.1  & (~\encrypt_mode<0>  & \encrypt<0> )) | (\$$COND520<0>0.1  & (\encrypt_mode<0>  & ~\encrypt<0> )),
  \[693]  = (\[672]  & (~\[524]  & ~\main_1/preS<14>0.1 )) | (\[623]  & \[530] ),
  \main_1/preS<34>0.1  = (~\data<55>  & \D<4> ) | (\data<55>  & ~\D<4> ),
  \$$COND359<0>376.1  = \[705]  & \[643] ,
  \$$COND249<0>226.1  = \[675]  & (\[627]  & ~\main_1/preS<19>0.1 ),
  \$$COND207<0>226.1  = \[669]  & \[664] ,
  \main_1/S1_1/$S1<2>76.1  = (~\[657]  & (~\[647]  & (~\[629]  & (~\[544]  & (~\[538]  & \main_1/preS<8>0.1 ))))) | ((~\[717]  & (~\[622]  & (\[523]  & (~\main_1/preS<8>0.1  & ~\main_1/preS<11>0.1 )))) | ((~\[647]  & (~\[646]  & (\[568]  & (~\[523]  & \main_1/preS<11>0.1 )))) | ((~\[717]  & (\[647]  & (~\[640]  & ~\[568] ))) | ((~\[717]  & (\[646]  & (\[523]  & ~\main_1/preS<8>0.1 ))) | ((~\[717]  & (~\[570]  & (\[538]  & \[523] ))) | ((\[717]  & (~\[515]  & (\main_1/preS<7>0.1  & \main_1/preS<11>0.1 ))) | ((~\[657]  & (~\[629]  & (\[622]  & ~\main_1/preS<11>0.1 ))) | (\[717]  & (\[544]  & ~\[508] ))))))))),
  \main_1/S7_1/$S7<2>526.1  = (~\[730]  & (~\[711]  & (~\[655]  & (~\[580]  & (~\[564]  & (~\[534]  & \main_1/preS<45>0.1 )))))) | ((~\[723]  & (\[583]  & (~\[560]  & \main_1/preS<44>0.1 ))) | ((~\[721]  & (~\[583]  & (\[560]  & ~\main_1/preS<46>0.1 ))) | ((~\[655]  & (~\[564]  & (\[549]  & \[517] ))) | ((\[723]  & (\[511]  & ~\main_1/preS<45>0.1 )) | ((\[652]  & (~\[517]  & ~\main_1/preS<45>0.1 )) | ((\[580]  & (\[513]  & \[511] )) | ((\[564]  & (\[560]  & ~\main_1/preS<45>0.1 )) | ((\[721]  & \[580] ) | (\[621]  & \[583] ))))))))),
  \$$COND40<0>1.1  = 0,
  \main_1/preS<47>0.1  = (~\data<32>  & \D<3> ) | (\data<32>  & ~\D<3> ),
  \main_1/preS<4>0.1  = (~\data<35>  & \C<0> ) | (\data<35>  & ~\C<0> ),
  \main_1/preS<30>0.1  = (~\data<51>  & \D<1> ) | (\data<51>  & ~\D<1> ),
  \main_1/S3_1/$S3<2>226.1  = (\[529]  & (\[510]  & (\main_1/preS<21>0.1  & ~\main_1/preS<20>0.1 ))) | ((~\[510]  & (\main_1/preS<23>0.1  & (~\main_1/preS<21>0.1  & \main_1/preS<20>0.1 ))) | ((\[664]  & (~\$$COND207<0>226.1  & ~\main_1/preS<23>0.1 )) | ((\[653]  & (\main_1/preS<23>0.1  & \main_1/preS<19>0.1 )) | ((\[641]  & (\main_1/preS<21>0.1  & \main_1/preS<19>0.1 )) | ((\[637]  & (~\$$COND232<0>226.1  & ~\main_1/preS<21>0.1 )) | ((\[628]  & (\[533]  & ~\$$COND232<0>226.1 )) | ((\[726]  & ~\main_1/preS<18>0.1 ) | ((\[704]  & \[627] ) | ((\[669]  & ~\[510] ) | ((\[650]  & \[535] ) | ((\[618]  & \[572] ) | (\$$COND258<0>226.1  | (\$$COND249<0>226.1  | (\$$COND225<0>226.1  | \$$COND216<0>226.1 )))))))))))))),
  \[10]  = (\[493]  & \inreg<38> ) | (\[492]  & \inreg<46> ),
  \[11]  = (\[493]  & \inreg<37> ) | (\[492]  & \inreg<45> ),
  \[12]  = (\[493]  & \inreg<36> ) | (\[492]  & \inreg<44> ),
  \[13]  = (\[493]  & \inreg<35> ) | (\[492]  & \inreg<43> ),
  \[14]  = (\[493]  & \inreg<34> ) | (\[492]  & \inreg<42> ),
  \[15]  = (\[493]  & \inreg<33> ) | (\[492]  & \inreg<41> ),
  \main_1/preS<43>0.1  = (~\data<60>  & \D<13> ) | (\data<60>  & ~\D<13> ),
  \[16]  = (\[493]  & \inreg<32> ) | (\[492]  & \inreg<40> ),
  \main_1/preS<0>0.1  = (~\data<63>  & \C<13> ) | (\data<63>  & ~\C<13> ),
  \[17]  = (\[493]  & \inreg<31> ) | (\[492]  & \inreg<39> ),
  \[18]  = (\[493]  & \inreg<30> ) | (\[492]  & \inreg<38> ),
  \[19]  = (\[493]  & \inreg<29> ) | (\[492]  & \inreg<37> ),
  \[20]  = (\[493]  & \inreg<28> ) | (\[492]  & \inreg<36> ),
  \[21]  = (\[493]  & \inreg<27> ) | (\[492]  & \inreg<35> ),
  \[22]  = (\[493]  & \inreg<26> ) | (\[492]  & \inreg<34> ),
  \[23]  = (\[493]  & \inreg<25> ) | (\[492]  & \inreg<33> ),
  \[24]  = (\[493]  & \inreg<24> ) | (\[492]  & \inreg<32> ),
  \[25]  = (\[493]  & \inreg<23> ) | (\[492]  & \inreg<31> ),
  \[26]  = (\[493]  & \inreg<22> ) | (\[492]  & \inreg<30> ),
  \[27]  = (\[493]  & \inreg<21> ) | (\[492]  & \inreg<29> ),
  \[28]  = (\[493]  & \inreg<20> ) | (\[492]  & \inreg<28> ),
  \main_1/preS<16>0.1  = (~\data<43>  & \C<25> ) | (\data<43>  & ~\C<25> ),
  \[100]  = (\[493]  & \outreg<28> ) | ((\[492]  & \outreg<20> ) | (\$$COND520<0>0.1  & \data<53> )),
  \[29]  = (\[493]  & \inreg<19> ) | (\[492]  & \inreg<27> ),
  \[101]  = (\[607]  & \$$COND520<0>0.1 ) | ((\[493]  & \outreg<27> ) | (\[492]  & \outreg<19> )),
  \[102]  = (\[493]  & \outreg<26> ) | ((\[492]  & \outreg<18> ) | (\$$COND520<0>0.1  & \data<45> )),
  \[103]  = (\[608]  & \$$COND520<0>0.1 ) | ((\[493]  & \outreg<25> ) | (\[492]  & \outreg<17> )),
  \[104]  = (\[493]  & \outreg<24> ) | ((\[492]  & \outreg<16> ) | (\$$COND520<0>0.1  & \data<37> )),
  \main_1/S2_1/$S2<0>151.1  = (\[558]  & (~\[507]  & (\main_1/preS<17>0.1  & \main_1/S2_1/$S2<1>151.1 ))) | ((\[558]  & (\main_1/preS<16>0.1  & (\main_1/preS<12>0.1  & ~\main_1/S2_1/$S2<1>151.1 ))) | ((~\[555]  & (\[547]  & (\[524]  & ~\[507] ))) | ((~\[530]  & (\[519]  & (\[507]  & \main_1/preS<16>0.1 ))) | ((\[530]  & (\[507]  & (\main_1/preS<14>0.1  & \main_1/S2_1/$S2<1>151.1 ))) | ((\[656]  & (\[555]  & ~\main_1/preS<16>0.1 )) | ((\[584]  & (~\[555]  & ~\[509] )) | ((\[582]  & (~\[519]  & ~\main_1/preS<16>0.1 )) | ((\[558]  & (~\main_1/preS<17>0.1  & ~\main_1/preS<16>0.1 )) | ((~\[519]  & (~\[509]  & \main_1/S2_1/$S2<1>151.1 )) | \$$COND180<0>151.1 ))))))))),
  \[105]  = (\[609]  & \$$COND520<0>0.1 ) | ((\[493]  & \outreg<23> ) | (\[492]  & \outreg<15> )),
  \[106]  = (\[493]  & \outreg<22> ) | ((\[492]  & \outreg<14> ) | (\$$COND520<0>0.1  & \data<62> )),
  \[107]  = (\[610]  & \$$COND520<0>0.1 ) | ((\[493]  & \outreg<21> ) | (\[492]  & \outreg<13> )),
  \[30]  = (\[493]  & \inreg<18> ) | (\[492]  & \inreg<26> ),
  \main_1/S5_1/$S5<3>376.1  = (~\[625]  & (\[525]  & (\main_1/preS<35>0.1  & \main_1/preS<30>0.1 ))) | ((\[636]  & (~\[505]  & \main_1/preS<31>0.1 )) | ((\[632]  & (\[539]  & ~\main_1/preS<34>0.1 )) | ((\[620]  & (\[531]  & ~\main_1/preS<32>0.1 )) | ((\[619]  & (~\[505]  & \main_1/preS<33>0.1 )) | ((\[545]  & (~\main_1/preS<32>0.1  & ~\main_1/preS<31>0.1 )) | ((\[539]  & (~\[505]  & ~\main_1/preS<33>0.1 )) | ((\[532]  & (~\[516]  & \main_1/preS<35>0.1 )) | ((\[702]  & \[578] ) | ((\[701]  & ~\main_1/preS<30>0.1 ) | ((\[670]  & \[525] ) | ((\[636]  & \[632] ) | ((\[635]  & ~\[516] ) | ((\[632]  & \[578] ) | ((\[625]  & ~\main_1/preS<33>0.1 ) | \$$COND358<0>376.1 )))))))))))))),
  \[108]  = (\[493]  & \outreg<20> ) | ((\[492]  & \outreg<12> ) | (\$$COND520<0>0.1  & \data<54> )),
  \[31]  = (\[493]  & \inreg<17> ) | (\[492]  & \inreg<25> ),
  \[109]  = (\[611]  & \$$COND520<0>0.1 ) | ((\[493]  & \outreg<19> ) | (\[492]  & \outreg<11> )),
  \[32]  = (\[493]  & \inreg<16> ) | (\[492]  & \inreg<24> ),
  \[33]  = (\[493]  & \inreg<15> ) | (\[492]  & \inreg<23> ),
  \[34]  = (\[493]  & \inreg<14> ) | (\[492]  & \inreg<22> ),
  \[35]  = (\[493]  & \inreg<13> ) | (\[492]  & \inreg<21> ),
  \[36]  = (\[493]  & \inreg<12> ) | (\[492]  & \inreg<20> ),
  \[37]  = (\[493]  & \inreg<11> ) | (\[492]  & \inreg<19> ),
  \main_1/S7_1/$S7<1>526.1  = (\[723]  & (\main_1/preS<45>0.1  & \main_1/S7_1/$S7<2>526.1 )) | ((\[655]  & (~\[559]  & \[549] )) | ((\[564]  & (\main_1/preS<47>0.1  & ~\main_1/S7_1/$S7<2>526.1 )) | ((~\[517]  & (~\main_1/preS<45>0.1  & ~\main_1/preS<43>0.1 )) | ((~\[511]  & (~\main_1/preS<43>0.1  & ~\main_1/preS<42>0.1 )) | ((\[731]  & ~\main_1/preS<44>0.1 ) | ((\[730]  & \main_1/preS<44>0.1 ) | ((\[721]  & \main_1/preS<43>0.1 ) | ((\[665]  & \[559] ) | ((\[649]  & \main_1/preS<45>0.1 ) | ((\[621]  & \[559] ) | (\[718]  | \$$COND484<0>526.1 ))))))))))),
  \[38]  = (\[493]  & \inreg<10> ) | (\[492]  & \inreg<18> ),
  \[110]  = (\[493]  & \outreg<18> ) | ((\[492]  & \outreg<10> ) | (\$$COND520<0>0.1  & \data<46> )),
  \[39]  = (\[493]  & \inreg<9> ) | (\[492]  & \inreg<17> ),
  \[111]  = (\[612]  & \$$COND520<0>0.1 ) | ((\[493]  & \outreg<17> ) | (\[492]  & \outreg<9> )),
  \main_1/preS<29>0.1  = (~\data<52>  & \D<26> ) | (\data<52>  & ~\D<26> ),
  \[112]  = (\[493]  & \outreg<16> ) | ((\[492]  & \outreg<8> ) | (\$$COND520<0>0.1  & \data<38> )),
  \[113]  = (\[613]  & \$$COND520<0>0.1 ) | ((\[493]  & \outreg<15> ) | (\[492]  & \outreg<7> )),
  \[114]  = (\[493]  & \outreg<14> ) | ((\[492]  & \outreg<6> ) | (\$$COND520<0>0.1  & \data<63> )),
  \[115]  = (\[614]  & \$$COND520<0>0.1 ) | ((\[493]  & \outreg<13> ) | (\[492]  & \outreg<5> )),
  \main_1/preS<12>0.1  = (~\data<39>  & \C<22> ) | (\data<39>  & ~\C<22> ),
  \[116]  = (\[493]  & \outreg<12> ) | ((\[492]  & \outreg<4> ) | (\$$COND520<0>0.1  & \data<55> )),
  \[117]  = (\[615]  & \$$COND520<0>0.1 ) | ((\[493]  & \outreg<11> ) | (\[492]  & \outreg<3> )),
  \[40]  = (\[493]  & \inreg<8> ) | (\[492]  & \inreg<16> ),
  \[118]  = (\[493]  & \outreg<10> ) | ((\[492]  & \outreg<2> ) | (\$$COND520<0>0.1  & \data<47> )),
  \[41]  = (\[493]  & \inreg<7> ) | (\[492]  & \inreg<15> ),
  \$$COND445<0>451.1  = \[633]  & (\[573]  & \main_1/preS<41>0.1 ),
  \[119]  = (\[616]  & \$$COND520<0>0.1 ) | ((\[493]  & \outreg<9> ) | (\[492]  & \outreg<1> )),
  \[42]  = (\[493]  & \inreg<6> ) | (\[492]  & \inreg<14> ),
  \main_1/preS<8>0.1  = (~\data<37>  & \C<14> ) | (\data<37>  & ~\C<14> ),
  \[43]  = (\[493]  & \inreg<5> ) | (\[492]  & \inreg<13> ),
  \[44]  = (\[493]  & \inreg<4> ) | (\[492]  & \inreg<12> ),
  \[45]  = (\[493]  & \inreg<3> ) | (\[492]  & \inreg<11> ),
  \[46]  = (\[493]  & \inreg<2> ) | (\[492]  & \inreg<10> ),
  \$$COND477<0>526.1  = \[711]  & \[580] ,
  \[47]  = (\[493]  & \inreg<1> ) | (\[492]  & \inreg<9> ),
  \[48]  = (\[493]  & \inreg<0> ) | (\[492]  & \inreg<8> ),
  \[120]  = (\[493]  & \outreg<8> ) | ((\[492]  & \outreg<0> ) | (\$$COND520<0>0.1  & \data<39> )),
  \[49]  = (\[493]  & \data_in<7> ) | (\[492]  & \inreg<7> ),
  \[500]  = \[495]  & ~\generate_key_1/shift_by_one<0>605.1 ,
  \[121]  = (\[613]  & ~\$$COND520<0>0.1 ) | (\$$COND520<0>0.1  & \data_in<6> ),
  \[501]  = \[496]  & ~\generate_key_1/shift_by_one<0>605.1 ,
  \[122]  = (\[609]  & ~\$$COND520<0>0.1 ) | (\$$COND520<0>0.1  & \inreg<6> ),
  \[502]  = \[496]  & \generate_key_1/shift_by_one<0>605.1 ,
  \[123]  = (\[605]  & ~\$$COND520<0>0.1 ) | (\$$COND520<0>0.1  & \inreg<14> ),
  \[503]  = \[495]  & \generate_key_1/shift_by_one<0>605.1 ,
  \[124]  = (\[601]  & ~\$$COND520<0>0.1 ) | (\$$COND520<0>0.1  & \inreg<22> ),
  \[504]  = \[630]  | \[581] ,
  \[125]  = (\[597]  & ~\$$COND520<0>0.1 ) | (\$$COND520<0>0.1  & \inreg<30> ),
  \[505]  = \main_1/preS<32>0.1  | \main_1/preS<30>0.1 ,
  \[126]  = (\[593]  & ~\$$COND520<0>0.1 ) | (\$$COND520<0>0.1  & \inreg<38> ),
  \main_1/S3_1/$S3<1>226.1  = (\[729]  & (\main_1/preS<22>0.1  & \main_1/preS<20>0.1 )) | ((\[653]  & (\main_1/preS<22>0.1  & \main_1/preS<19>0.1 )) | ((\[641]  & (\[628]  & ~\main_1/preS<21>0.1 )) | ((\[627]  & (\[551]  & \main_1/preS<19>0.1 )) | ((\[618]  & (\[529]  & ~\main_1/preS<19>0.1 )) | ((\[618]  & (~\main_1/preS<21>0.1  & ~\main_1/preS<19>0.1 )) | ((\[535]  & (\[533]  & ~\$$COND196<0>226.1 )) | ((\[726]  & \main_1/preS<20>0.1 ) | ((\[712]  & \main_1/preS<19>0.1 ) | ((\[654]  & \[627] ) | ((\[651]  & \[579] ) | (\$$COND254<0>226.1  | (\$$COND207<0>226.1  | (\$$COND258<0>226.1  | (\$$COND238<0>226.1  | (\$$COND233<0>226.1  | \$$COND210<0>226.1 ))))))))))))))),
  \[506]  = \[575]  | \[556] ,
  \[127]  = (\[589]  & ~\$$COND520<0>0.1 ) | (\$$COND520<0>0.1  & \inreg<46> ),
  \[50]  = (\[493]  & \data_in<6> ) | (\[492]  & \inreg<6> ),
  \[507]  = (\main_1/preS<14>0.1  & ~\main_1/preS<13>0.1 ) | \[707] ,
  \main_1/preS<25>0.1  = (~\data<48>  & \D<23> ) | (\data<48>  & ~\D<23> ),
  \[128]  = (\[585]  & ~\$$COND520<0>0.1 ) | (\$$COND520<0>0.1  & \inreg<54> ),
  \[51]  = (\[493]  & \data_in<5> ) | (\[492]  & \inreg<5> ),
  \[508]  = ~\main_1/preS<9>0.1  | ~\main_1/preS<7>0.1 ,
  \$$COND210<0>226.1  = \[641]  & (\[626]  & \[551] ),
  \main_1/S6_1/$S6<3>451.1  = (\[645]  & (\main_1/preS<39>0.1  & (\main_1/preS<37>0.1  & ~\main_1/S6_1/$S6<2>451.1 ))) | ((\[550]  & (~\main_1/preS<39>0.1  & (\main_1/preS<38>0.1  & \main_1/S6_1/$S6<2>451.1 ))) | ((\main_1/preS<40>0.1  & (~\main_1/preS<38>0.1  & (\main_1/preS<36>0.1  & ~\main_1/S6_1/$S6<2>451.1 ))) | ((\[667]  & (\[644]  & ~\main_1/preS<40>0.1 )) | ((\[722]  & ~\[639] ) | ((\[722]  & ~\[573] ) | ((\[719]  & ~\main_1/preS<37>0.1 ) | ((\[713]  & ~\main_1/preS<37>0.1 ) | ((\[639]  & ~\main_1/S6_1/$S6<2>451.1 ) | ((\[634]  & ~\main_1/preS<36>0.1 ) | ((\[633]  & \[550] ) | ((\[631]  & \[577] ) | (\[682]  | \$$COND414<0>451.1 )))))))))))),
  \[129]  = (\[614]  & ~\$$COND520<0>0.1 ) | (\$$COND520<0>0.1  & \data_in<4> ),
  \[52]  = (\[493]  & \data_in<4> ) | (\[492]  & \inreg<4> ),
  \[509]  = \main_1/preS<15>0.1  | \main_1/preS<13>0.1 ,
  \[53]  = (\[493]  & \data_in<3> ) | (\[492]  & \inreg<3> ),
  \main_1/S0_1/$S0<1>1.1  = (~\[566]  & (~\[557]  & (~\[548]  & (~\[537]  & \[536] )))) | ((\[567]  & (\[562]  & (~\[536]  & ~\[520] ))) | ((~\[557]  & (~\[537]  & (~\[528]  & \[518] ))) | ((\[709]  & (~\[561]  & \[528] )) | ((\[566]  & (\[557]  & \[528] )) | ((\[561]  & (\[548]  & \[537] )) | ((\[557]  & (\[548]  & \[536] )) | ((\[557]  & (~\[528]  & ~\[518] )) | ((\[714]  & \main_1/preS<4>0.1 ) | ((\[706]  & \[554] ) | ((\[677]  & \[566] ) | (~\[562]  & \[548] ))))))))))),
  \[54]  = (\[493]  & \data_in<2> ) | (\[492]  & \inreg<2> ),
  \[55]  = (\[493]  & \data_in<1> ) | (\[492]  & \inreg<1> ),
  \[56]  = (\[493]  & \data_in<0> ) | (\[492]  & \inreg<0> ),
  \inreg_new<50>  = \[6] ,
  \[57]  = (\[585]  & \$$COND520<0>0.1 ) | (\[492]  & \outreg<63> ),
  \[58]  = (\[492]  & \outreg<62> ) | (\$$COND520<0>0.1  & \data<56> ),
  \main_1/preS<37>0.1  = (~\data<56>  & \D<20> ) | (\data<56>  & ~\D<20> ),
  \[130]  = (\[610]  & ~\$$COND520<0>0.1 ) | (\$$COND520<0>0.1  & \inreg<4> ),
  \[59]  = (\[586]  & \$$COND520<0>0.1 ) | (\[492]  & \outreg<61> ),
  \[510]  = ~\main_1/preS<19>0.1  | ~\main_1/preS<18>0.1 ,
  \inreg_new<9>  = \[47] ,
  \[131]  = (\[606]  & ~\$$COND520<0>0.1 ) | (\$$COND520<0>0.1  & \inreg<12> ),
  \[511]  = \main_1/preS<46>0.1  | ~\main_1/preS<44>0.1 ,
  \[701]  = \[620]  & ~\main_1/preS<31>0.1 ,
  \inreg_new<54>  = \[2] ,
  \[132]  = (\[602]  & ~\$$COND520<0>0.1 ) | (\$$COND520<0>0.1  & \inreg<20> ),
  \[512]  = \main_1/preS<39>0.1  & \main_1/preS<36>0.1 ,
  \[702]  = \[539]  & \main_1/preS<32>0.1 ,
  \inreg_new<53>  = \[3] ,
  \[133]  = (\[598]  & ~\$$COND520<0>0.1 ) | (\$$COND520<0>0.1  & \inreg<28> ),
  \[513]  = \main_1/preS<45>0.1  & \main_1/preS<42>0.1 ,
  \[703]  = \[553]  & \main_1/preS<28>0.1 ,
  \inreg_new<52>  = \[4] ,
  \inreg_new<6>  = \[50] ,
  \[134]  = (\[594]  & ~\$$COND520<0>0.1 ) | (\$$COND520<0>0.1  & \inreg<36> ),
  \[514]  = ~\main_1/preS<40>0.1  | \main_1/preS<39>0.1 ,
  \[704]  = \[579]  & \main_1/preS<21>0.1 ,
  \inreg_new<51>  = \[5] ,
  \inreg_new<5>  = \[51] ,
  \[135]  = (\[590]  & ~\$$COND520<0>0.1 ) | (\$$COND520<0>0.1  & \inreg<44> ),
  \[515]  = \main_1/preS<8>0.1  | ~\main_1/preS<6>0.1 ,
  \[705]  = \[671]  & ~\main_1/preS<31>0.1 ,
  \inreg_new<8>  = \[48] ,
  \[136]  = (\[586]  & ~\$$COND520<0>0.1 ) | (\$$COND520<0>0.1  & \inreg<52> ),
  \[516]  = ~\main_1/preS<32>0.1  | \main_1/preS<30>0.1 ,
  \[706]  = ~\[518]  & \main_1/preS<2>0.1 ,
  \inreg_new<7>  = \[49] ,
  \[137]  = (\[615]  & ~\$$COND520<0>0.1 ) | (\$$COND520<0>0.1  & \data_in<2> ),
  \[60]  = (\[492]  & \outreg<60> ) | (\$$COND520<0>0.1  & \data<48> ),
  \[517]  = ~\main_1/preS<46>0.1  | \main_1/preS<42>0.1 ,
  \[707]  = ~\main_1/preS<14>0.1  & \main_1/preS<13>0.1 ,
  \inreg_new<2>  = \[54] ,
  \[138]  = (\[611]  & ~\$$COND520<0>0.1 ) | (\$$COND520<0>0.1  & \inreg<2> ),
  \[61]  = (\[587]  & \$$COND520<0>0.1 ) | (\[492]  & \outreg<59> ),
  \[518]  = ~\main_1/preS<3>0.1  | \main_1/preS<1>0.1 ,
  \inreg_new<55>  = \[1] ,
  \inreg_new<1>  = \[55] ,
  \[139]  = (\[607]  & ~\$$COND520<0>0.1 ) | (\$$COND520<0>0.1  & \inreg<10> ),
  \[62]  = (\[492]  & \outreg<58> ) | (\$$COND520<0>0.1  & \data<40> ),
  \$$COND317<0>301.1  = 0,
  \[519]  = ~\main_1/preS<17>0.1  | \main_1/preS<12>0.1 ,
  \[709]  = \[566]  & \[537] ,
  \inreg_new<4>  = \[52] ,
  \[63]  = (\[588]  & \$$COND520<0>0.1 ) | (\[492]  & \outreg<57> ),
  \inreg_new<3>  = \[53] ,
  \[64]  = (\[492]  & \outreg<56> ) | (\$$COND520<0>0.1  & \data<32> ),
  \[65]  = (\[589]  & \$$COND520<0>0.1 ) | ((\[493]  & \outreg<63> ) | (\[492]  & \outreg<55> )),
  \[66]  = (\[493]  & \outreg<62> ) | ((\[492]  & \outreg<54> ) | (\$$COND520<0>0.1  & \data<57> )),
  \inreg_new<0>  = \[56] ,
  \[67]  = (\[590]  & \$$COND520<0>0.1 ) | ((\[493]  & \outreg<61> ) | (\[492]  & \outreg<53> )),
  \main_1/preS<21>0.1  = (~\data<46>  & \C<19> ) | (\data<46>  & ~\C<19> ),
  \[68]  = (\[493]  & \outreg<60> ) | ((\[492]  & \outreg<52> ) | (\$$COND520<0>0.1  & \data<49> )),
  \[140]  = (\[603]  & ~\$$COND520<0>0.1 ) | (\$$COND520<0>0.1  & \inreg<18> ),
  \[69]  = (\[591]  & \$$COND520<0>0.1 ) | ((\[493]  & \outreg<59> ) | (\[492]  & \outreg<51> )),
  \[520]  = \main_1/preS<5>0.1  & \main_1/preS<4>0.1 ,
  \[710]  = \[568]  & \main_1/preS<10>0.1 ,
  \[141]  = (\[599]  & ~\$$COND520<0>0.1 ) | (\$$COND520<0>0.1  & \inreg<26> ),
  \generate_key_1/shift_by_one<0>605.1  = (~\[648]  & (~\count<1>  & ~\count<2> )) | (\[648]  & (\count<1>  & \count<2> )),
  \[521]  = \main_1/preS<26>0.1  & ~\main_1/preS<25>0.1 ,
  \[711]  = \[583]  & ~\[511] ,
  \[142]  = (\[595]  & ~\$$COND520<0>0.1 ) | (\$$COND520<0>0.1  & \inreg<34> ),
  \[522]  = \main_1/preS<38>0.1  | \main_1/preS<37>0.1 ,
  \[712]  = \[572]  & \main_1/preS<20>0.1 ,
  \[143]  = (\[591]  & ~\$$COND520<0>0.1 ) | (\$$COND520<0>0.1  & \inreg<42> ),
  \[523]  = \main_1/preS<6>0.1  | \main_1/preS<10>0.1 ,
  \[713]  = \[574]  & \[512] ,
  \[144]  = (\[587]  & ~\$$COND520<0>0.1 ) | (\$$COND520<0>0.1  & \inreg<50> ),
  \[524]  = ~\main_1/preS<17>0.1  | ~\main_1/preS<12>0.1 ,
  \[714]  = \[561]  & ~\[518] ,
  \[145]  = (\[616]  & ~\$$COND520<0>0.1 ) | (\$$COND520<0>0.1  & \data_in<0> ),
  \[525]  = \main_1/preS<34>0.1  & \main_1/preS<33>0.1 ,
  \main_1/preS<33>0.1  = (~\data<54>  & \D<16> ) | (\data<54>  & ~\D<16> ),
  \[715]  = \[584]  & ~\[524] ,
  \[146]  = (\[612]  & ~\$$COND520<0>0.1 ) | (\$$COND520<0>0.1  & \inreg<0> ),
  \$$COND286<0>301.1  = 0,
  \[526]  = ~\main_1/preS<28>0.1  & ~\main_1/preS<24>0.1 ,
  \[716]  = \[633]  & ~\main_1/preS<41>0.1 ,
  \[147]  = (\[608]  & ~\$$COND520<0>0.1 ) | (\$$COND520<0>0.1  & \inreg<8> ),
  \[70]  = (\[493]  & \outreg<58> ) | ((\[492]  & \outreg<50> ) | (\$$COND520<0>0.1  & \data<41> )),
  \[527]  = ~\main_1/preS<28>0.1  | ~\main_1/preS<24>0.1 ,
  \[717]  = \main_1/preS<6>0.1  & \main_1/preS<10>0.1 ,
  \[148]  = (\[604]  & ~\$$COND520<0>0.1 ) | (\$$COND520<0>0.1  & \inreg<16> ),
  \[71]  = (\[592]  & \$$COND520<0>0.1 ) | ((\[493]  & \outreg<57> ) | (\[492]  & \outreg<49> )),
  \$$COND254<0>226.1  = \[704]  & \[529] ,
  \[528]  = \main_1/preS<2>0.1  | \main_1/preS<0>0.1 ,
  \[718]  = \[652]  & \[513] ,
  \encrypt_mode_new<0>  = \[245] ,
  \[149]  = (\[600]  & ~\$$COND520<0>0.1 ) | (\$$COND520<0>0.1  & \inreg<24> ),
  \[72]  = (\[493]  & \outreg<56> ) | ((\[492]  & \outreg<48> ) | (\$$COND520<0>0.1  & \data<33> )),
  \[529]  = \main_1/preS<23>0.1  & \main_1/preS<22>0.1 ,
  \[719]  = \[577]  & ~\main_1/preS<41>0.1 ,
  \[73]  = (\[593]  & \$$COND520<0>0.1 ) | ((\[493]  & \outreg<55> ) | (\[492]  & \outreg<47> )),
  \[74]  = (\[493]  & \outreg<54> ) | ((\[492]  & \outreg<46> ) | (\$$COND520<0>0.1  & \data<58> )),
  \[75]  = (\[594]  & \$$COND520<0>0.1 ) | ((\[493]  & \outreg<53> ) | (\[492]  & \outreg<45> )),
  \outreg_new<9>  = \[111] ,
  \[76]  = (\[493]  & \outreg<52> ) | ((\[492]  & \outreg<44> ) | (\$$COND520<0>0.1  & \data<50> )),
  \[77]  = (\[595]  & \$$COND520<0>0.1 ) | ((\[493]  & \outreg<51> ) | (\[492]  & \outreg<43> )),
  \outreg_new<51>  = \[69] ,
  \[78]  = (\[493]  & \outreg<50> ) | ((\[492]  & \outreg<42> ) | (\$$COND520<0>0.1  & \data<42> )),
  \outreg_new<52>  = \[68] ,
  \[150]  = (\[596]  & ~\$$COND520<0>0.1 ) | (\$$COND520<0>0.1  & \inreg<32> ),
  \[79]  = (\[596]  & \$$COND520<0>0.1 ) | ((\[493]  & \outreg<49> ) | (\[492]  & \outreg<41> )),
  \outreg_new<53>  = \[67] ,
  \[530]  = ~\main_1/preS<17>0.1  & \main_1/preS<12>0.1 ,
  \outreg_new<5>  = \[115] ,
  \[720]  = \[624]  & ~\[514] ,
  \[151]  = (\[592]  & ~\$$COND520<0>0.1 ) | (\$$COND520<0>0.1  & \inreg<40> ),
  \outreg_new<54>  = \[66] ,
  \[531]  = \main_1/preS<31>0.1  & \main_1/preS<30>0.1 ,
  \outreg_new<6>  = \[114] ,
  \[721]  = \[559]  & ~\[511] ,
  \[152]  = (\[588]  & ~\$$COND520<0>0.1 ) | (\$$COND520<0>0.1  & \inreg<48> ),
  \[532]  = \main_1/preS<34>0.1  & ~\main_1/preS<33>0.1 ,
  \outreg_new<7>  = \[113] ,
  \[722]  = \[573]  & \[542] ,
  \main_1/S4_1/$S4<0>301.1  = (~\[660]  & (~\[565]  & (~\[553]  & (\[506]  & ~\main_1/preS<25>0.1 )))) | ((~\[725]  & (\[576]  & (~\[553]  & \main_1/preS<28>0.1 ))) | ((\[630]  & (~\[565]  & (\[556]  & ~\[553] ))) | ((\[630]  & (\[553]  & \main_1/preS<24>0.1 )) | ((\[581]  & (\[540]  & \main_1/preS<28>0.1 )) | ((\[576]  & (\[575]  & \[565] )) | ((\[565]  & (~\[506]  & \main_1/preS<26>0.1 )) | ((\[526]  & (~\[504]  & \main_1/preS<27>0.1 )) | ((\[728]  & \[546] ) | ((\[703]  & ~\[527] ) | (\[703]  & \[521] )))))))))),
  \[153]  = (\data_in<7>  & \$$COND520<0>0.1 ) | (\data<63>  & ~\$$COND520<0>0.1 ),
  \[533]  = ~\main_1/preS<23>0.1  & ~\main_1/preS<19>0.1 ,
  \outreg_new<8>  = \[112] ,
  \[723]  = \main_1/preS<47>0.1  & \main_1/preS<43>0.1 ,
  \[154]  = (\inreg<7>  & \$$COND520<0>0.1 ) | (\data<62>  & ~\$$COND520<0>0.1 ),
  \[534]  = \main_1/preS<47>0.1  & ~\main_1/preS<44>0.1 ,
  \outreg_new<1>  = \[119] ,
  \[724]  = \[571]  & ~\[508] ,
  \[155]  = (\inreg<15>  & \$$COND520<0>0.1 ) | (\data<61>  & ~\$$COND520<0>0.1 ),
  \outreg_new<50>  = \[70] ,
  \[535]  = ~\main_1/preS<20>0.1  & ~\main_1/preS<18>0.1 ,
  \outreg_new<2>  = \[118] ,
  \[725]  = \[556]  & \[546] ,
  \[156]  = (\inreg<23>  & \$$COND520<0>0.1 ) | (\data<60>  & ~\$$COND520<0>0.1 ),
  \outreg_new<59>  = \[61] ,
  \[536]  = ~\main_1/preS<2>0.1  & \main_1/preS<0>0.1 ,
  \outreg_new<3>  = \[117] ,
  \[726]  = \[668]  & \[552] ,
  \[157]  = (\inreg<31>  & \$$COND520<0>0.1 ) | (\data<59>  & ~\$$COND520<0>0.1 ),
  \[80]  = (\[493]  & \outreg<48> ) | ((\[492]  & \outreg<40> ) | (\$$COND520<0>0.1  & \data<34> )),
  \[537]  = ~\main_1/preS<5>0.1  & \main_1/preS<4>0.1 ,
  \outreg_new<4>  = \[116] ,
  \[727]  = ~\[522]  & ~\main_1/preS<36>0.1 ,
  \main_1/preS<46>0.1  = (~\data<63>  & \D<0> ) | (\data<63>  & ~\D<0> ),
  \[158]  = (\inreg<39>  & \$$COND520<0>0.1 ) | (\data<58>  & ~\$$COND520<0>0.1 ),
  \[81]  = (\[597]  & \$$COND520<0>0.1 ) | ((\[493]  & \outreg<47> ) | (\[492]  & \outreg<39> )),
  \[538]  = \main_1/preS<9>0.1  & ~\main_1/preS<7>0.1 ,
  \[728]  = \[526]  & \main_1/preS<25>0.1 ,
  \$$COND232<0>226.1  = \[637]  & (\[628]  & ~\main_1/preS<21>0.1 ),
  \main_1/preS<3>0.1  = (~\data<34>  & \C<23> ) | (\data<34>  & ~\C<23> ),
  \[159]  = (\inreg<47>  & \$$COND520<0>0.1 ) | (\data<57>  & ~\$$COND520<0>0.1 ),
  \[82]  = (\[493]  & \outreg<46> ) | ((\[492]  & \outreg<38> ) | (\$$COND520<0>0.1  & \data<59> )),
  \[539]  = \main_1/preS<35>0.1  & ~\main_1/preS<31>0.1 ,
  \[729]  = ~\main_1/preS<19>0.1  & ~\main_1/preS<18>0.1 ,
  \[83]  = (\[598]  & \$$COND520<0>0.1 ) | ((\[493]  & \outreg<45> ) | (\[492]  & \outreg<37> )),
  \outreg_new<55>  = \[65] ,
  \data_new<43>  = \[141] ,
  \[84]  = (\[493]  & \outreg<44> ) | ((\[492]  & \outreg<36> ) | (\$$COND520<0>0.1  & \data<51> )),
  \outreg_new<56>  = \[64] ,
  \data_new<44>  = \[140] ,
  \outreg_new<0>  = \[120] ,
  \[85]  = (\[599]  & \$$COND520<0>0.1 ) | ((\[493]  & \outreg<43> ) | (\[492]  & \outreg<35> )),
  \outreg_new<57>  = \[63] ,
  \data_new<41>  = \[143] ,
  \[86]  = (\[493]  & \outreg<42> ) | ((\[492]  & \outreg<34> ) | (\$$COND520<0>0.1  & \data<43> )),
  \outreg_new<58>  = \[62] ,
  \data_new<42>  = \[142] ,
  \inreg_new<20>  = \[36] ,
  \[87]  = (\[600]  & \$$COND520<0>0.1 ) | ((\[493]  & \outreg<41> ) | (\[492]  & \outreg<33> )),
  \outreg_new<61>  = \[59] ,
  \[88]  = (\[493]  & \outreg<40> ) | ((\[492]  & \outreg<32> ) | (\$$COND520<0>0.1  & \data<35> )),
  \outreg_new<62>  = \[58] ,
  \data_new<40>  = \[144] ,
  \[160]  = (\inreg<55>  & \$$COND520<0>0.1 ) | (\data<56>  & ~\$$COND520<0>0.1 ),
  \main_1/S2_1/$S2<2>151.1  = (~\[672]  & (~\[663]  & (\[530]  & \main_1/preS<16>0.1 ))) | ((~\[623]  & (~\[617]  & (\[541]  & ~\[524] ))) | ((~\[623]  & (~\[584]  & (\[555]  & ~\main_1/preS<13>0.1 ))) | ((\[707]  & (\[582]  & ~\main_1/preS<12>0.1 )) | ((~\[617]  & (~\[541]  & ~\[519] )) | ((\[617]  & (~\[541]  & ~\[524] )) | ((\[541]  & (~\[519]  & ~\[509] )) | ((\[530]  & (~\[507]  & ~\main_1/preS<16>0.1 )) | (\[672]  & \[555] )))))))),
  \[89]  = (\[601]  & \$$COND520<0>0.1 ) | ((\[493]  & \outreg<39> ) | (\[492]  & \outreg<31> )),
  \outreg_new<63>  = \[57] ,
  \[540]  = ~\main_1/preS<29>0.1  & \main_1/preS<27>0.1 ,
  \[730]  = \[560]  & \[513] ,
  \[161]  = (\data_in<5>  & \$$COND520<0>0.1 ) | (\data<55>  & ~\$$COND520<0>0.1 ),
  \[541]  = \main_1/preS<16>0.1  | ~\main_1/preS<14>0.1 ,
  \[731]  = \[560]  & \[559] ,
  \inreg_new<24>  = \[32] ,
  \[162]  = (\inreg<5>  & \$$COND520<0>0.1 ) | (\data<54>  & ~\$$COND520<0>0.1 ),
  \[542]  = ~\main_1/preS<41>0.1  & ~\main_1/preS<40>0.1 ,
  \[732]  = \[544]  & \main_1/preS<8>0.1 ,
  \inreg_new<23>  = \[33] ,
  \[163]  = (\inreg<13>  & \$$COND520<0>0.1 ) | (\data<53>  & ~\$$COND520<0>0.1 ),
  \[543]  = ~\main_1/preS<9>0.1  & \main_1/preS<11>0.1 ,
  \inreg_new<22>  = \[34] ,
  \[164]  = (\inreg<21>  & \$$COND520<0>0.1 ) | (\data<52>  & ~\$$COND520<0>0.1 ),
  \[544]  = ~\main_1/preS<11>0.1  & \main_1/preS<10>0.1 ,
  \data_new<49>  = \[135] ,
  \inreg_new<21>  = \[35] ,
  \[165]  = (\inreg<29>  & \$$COND520<0>0.1 ) | (\data<51>  & ~\$$COND520<0>0.1 ),
  \outreg_new<60>  = \[60] ,
  \[545]  = ~\main_1/preS<35>0.1  & ~\main_1/preS<34>0.1 ,
  \inreg_new<28>  = \[28] ,
  \[166]  = (\inreg<37>  & \$$COND520<0>0.1 ) | (\data<50>  & ~\$$COND520<0>0.1 ),
  \[546]  = \main_1/preS<29>0.1  & ~\main_1/preS<27>0.1 ,
  \data_new<47>  = \[137] ,
  \inreg_new<27>  = \[29] ,
  \[167]  = (\inreg<45>  & \$$COND520<0>0.1 ) | (\data<49>  & ~\$$COND520<0>0.1 ),
  \[90]  = (\[493]  & \outreg<38> ) | ((\[492]  & \outreg<30> ) | (\$$COND520<0>0.1  & \data<60> )),
  \[547]  = \main_1/preS<16>0.1  & \main_1/preS<15>0.1 ,
  \data_new<48>  = \[136] ,
  \inreg_new<26>  = \[30] ,
  \[168]  = (\inreg<53>  & \$$COND520<0>0.1 ) | (\data<48>  & ~\$$COND520<0>0.1 ),
  \[91]  = (\[602]  & \$$COND520<0>0.1 ) | ((\[493]  & \outreg<37> ) | (\[492]  & \outreg<29> )),
  \[548]  = ~\main_1/preS<3>0.1  & ~\main_1/preS<1>0.1 ,
  \data_new<45>  = \[139] ,
  \inreg_new<25>  = \[31] ,
  \$$COND233<0>226.1  = \[675]  & \[650] ,
  \[169]  = (\data_in<3>  & \$$COND520<0>0.1 ) | (\data<47>  & ~\$$COND520<0>0.1 ),
  \[92]  = (\[493]  & \outreg<36> ) | ((\[492]  & \outreg<28> ) | (\$$COND520<0>0.1  & \data<52> )),
  \[549]  = ~\main_1/preS<47>0.1  & \main_1/preS<43>0.1 ,
  \data_new<46>  = \[138] ,
  \[93]  = (\[603]  & \$$COND520<0>0.1 ) | ((\[493]  & \outreg<35> ) | (\[492]  & \outreg<27> )),
  \data_new<33>  = \[151] ,
  \main_1/preS<19>0.1  = (~\data<44>  & \C<6> ) | (\data<44>  & ~\C<6> ),
  \[94]  = (\[493]  & \outreg<34> ) | ((\[492]  & \outreg<26> ) | (\$$COND520<0>0.1  & \data<44> )),
  \data_new<34>  = \[150] ,
  \[95]  = (\[604]  & \$$COND520<0>0.1 ) | ((\[493]  & \outreg<33> ) | (\[492]  & \outreg<25> )),
  \data_new<31>  = \[153] ,
  \inreg_new<29>  = \[27] ,
  \[96]  = (\[493]  & \outreg<32> ) | ((\[492]  & \outreg<24> ) | (\$$COND520<0>0.1  & \data<36> )),
  \data_new<32>  = \[152] ,
  \inreg_new<10>  = \[46] ,
  \[97]  = (\[605]  & \$$COND520<0>0.1 ) | ((\[493]  & \outreg<31> ) | (\[492]  & \outreg<23> )),
  \main_1/preS<42>0.1  = (~\data<59>  & \D<17> ) | (\data<59>  & ~\D<17> ),
  \[98]  = (\[493]  & \outreg<30> ) | ((\[492]  & \outreg<22> ) | (\$$COND520<0>0.1  & \data<61> )),
  \data_new<30>  = \[154] ,
  \[170]  = (\inreg<3>  & \$$COND520<0>0.1 ) | (\data<46>  & ~\$$COND520<0>0.1 ),
  \[99]  = (\[606]  & \$$COND520<0>0.1 ) | ((\[493]  & \outreg<29> ) | (\[492]  & \outreg<21> )),
  \[550]  = \main_1/preS<41>0.1  & \main_1/preS<37>0.1 ,
  \[171]  = (\inreg<11>  & \$$COND520<0>0.1 ) | (\data<45>  & ~\$$COND520<0>0.1 ),
  \[551]  = \main_1/preS<21>0.1  & \main_1/preS<20>0.1 ,
  \inreg_new<14>  = \[42] ,
  \[172]  = (\inreg<19>  & \$$COND520<0>0.1 ) | (\data<44>  & ~\$$COND520<0>0.1 ),
  \[552]  = ~\main_1/preS<22>0.1  & ~\main_1/preS<21>0.1 ,
  \inreg_new<13>  = \[43] ,
  \[173]  = (\inreg<27>  & \$$COND520<0>0.1 ) | (\data<43>  & ~\$$COND520<0>0.1 ),
  \[553]  = \main_1/preS<29>0.1  & \main_1/preS<27>0.1 ,
  \inreg_new<12>  = \[44] ,
  \[174]  = (\inreg<35>  & \$$COND520<0>0.1 ) | (\data<42>  & ~\$$COND520<0>0.1 ),
  \[554]  = ~\main_1/preS<5>0.1  & ~\main_1/preS<4>0.1 ,
  \data_new<39>  = \[145] ,
  \inreg_new<11>  = \[45] ,
  \[175]  = (\inreg<43>  & \$$COND520<0>0.1 ) | (\data<41>  & ~\$$COND520<0>0.1 ),
  \[555]  = ~\main_1/preS<17>0.1  & ~\main_1/preS<12>0.1 ,
  \inreg_new<18>  = \[38] ,
  \[176]  = (\inreg<51>  & \$$COND520<0>0.1 ) | (\data<40>  & ~\$$COND520<0>0.1 ),
  \[556]  = \main_1/preS<28>0.1  & ~\main_1/preS<24>0.1 ,
  \data_new<37>  = \[147] ,
  \inreg_new<17>  = \[39] ,
  \[177]  = (\data_in<1>  & \$$COND520<0>0.1 ) | (\data<39>  & ~\$$COND520<0>0.1 ),
  \[557]  = \main_1/preS<5>0.1  & ~\main_1/preS<4>0.1 ,
  \data_new<38>  = \[146] ,
  \inreg_new<16>  = \[40] ,
  \[178]  = (\inreg<1>  & \$$COND520<0>0.1 ) | (\data<38>  & ~\$$COND520<0>0.1 ),
  \[558]  = ~\main_1/preS<15>0.1  & \main_1/preS<13>0.1 ,
  \data_new<35>  = \[149] ,
  \inreg_new<15>  = \[41] ,
  \[179]  = (\inreg<9>  & \$$COND520<0>0.1 ) | (\data<37>  & ~\$$COND520<0>0.1 ),
  \[559]  = ~\main_1/preS<45>0.1  & \main_1/preS<42>0.1 ,
  \data_new<36>  = \[148] ,
  \data_new<23>  = \[161] ,
  \data_new<24>  = \[160] ,
  \data_new<21>  = \[163] ,
  \inreg_new<19>  = \[37] ,
  \data_new<22>  = \[162] ,
  \inreg_new<40>  = \[16] ,
  \data_new<20>  = \[164] ,
  \[180]  = (\inreg<17>  & \$$COND520<0>0.1 ) | (\data<36>  & ~\$$COND520<0>0.1 ),
  \[560]  = ~\main_1/preS<47>0.1  & ~\main_1/preS<43>0.1 ,
  \main_1/preS<15>0.1  = (~\data<42>  & \C<3> ) | (\data<42>  & ~\C<3> ),
  \[181]  = (\inreg<25>  & \$$COND520<0>0.1 ) | (\data<35>  & ~\$$COND520<0>0.1 ),
  \[561]  = \main_1/preS<2>0.1  & \main_1/preS<0>0.1 ,
  \inreg_new<44>  = \[12] ,
  \[182]  = (\inreg<33>  & \$$COND520<0>0.1 ) | (\data<34>  & ~\$$COND520<0>0.1 ),
  \[562]  = ~\main_1/preS<2>0.1  | \main_1/preS<0>0.1 ,
  \inreg_new<43>  = \[13] ,
  \[183]  = (\inreg<41>  & \$$COND520<0>0.1 ) | (\data<33>  & ~\$$COND520<0>0.1 ),
  \inreg_new<42>  = \[14] ,
  \[184]  = (\inreg<49>  & \$$COND520<0>0.1 ) | (\data<32>  & ~\$$COND520<0>0.1 ),
  \[564]  = \main_1/preS<46>0.1  & \main_1/preS<44>0.1 ,
  \data_new<29>  = \[155] ,
  \inreg_new<41>  = \[15] ,
  \[185]  = (\[490]  & (\generate_key_1/shift_by_one<0>605.1  & (~\$$COND520<0>0.1  & \count<1> ))) | (\[490]  & (~\generate_key_1/shift_by_one<0>605.1  & \count<3> )),
  \[565]  = ~\main_1/preS<29>0.1  & ~\main_1/preS<27>0.1 ,
  \inreg_new<48>  = \[8] ,
  \[186]  = (\[490]  & (~\[188]  & (\count<1>  & ~\count<2> ))) | ((\[188]  & \count<2> ) | (\[187]  & \count<2> )),
  \[566]  = \main_1/preS<3>0.1  & \main_1/preS<1>0.1 ,
  \data_new<27>  = \[157] ,
  \inreg_new<47>  = \[9] ,
  \[187]  = (\[490]  & (~\[188]  & ~\count<1> )) | (\[188]  & \count<1> ),
  \[567]  = ~\main_1/preS<3>0.1  & \main_1/preS<1>0.1 ,
  \data_new<28>  = \[156] ,
  \inreg_new<46>  = \[10] ,
  \[188]  = \[490]  & ~\count<0> ;
endmodule

