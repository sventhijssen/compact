// IWLS benchmark module "comp" printed on Wed May 29 16:07:21 2002
module comp(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, \x , y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0);
input
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  t,
  u,
  v,
  w,
  \x ,
  y,
  z,
  a0,
  b0,
  c0,
  d0,
  e0,
  f0;
output
  g0,
  h0,
  i0;
wire
  k1,
  k2,
  l1,
  l2,
  m0,
  m1,
  m2,
  n1,
  n2,
  o0,
  o1,
  o2,
  p1,
  p2,
  \[0] ,
  q0,
  q1,
  q2,
  \[1] ,
  r1,
  r2,
  \[2] ,
  s0,
  s1,
  s2,
  u0,
  v0,
  w0,
  x0,
  x1,
  x2,
  y0,
  y1,
  y2,
  z0,
  z1,
  z2,
  a1,
  a2,
  a3,
  b1,
  b2,
  b3,
  c1,
  c2,
  c3,
  d1,
  d2,
  d3,
  e1,
  e2,
  e3,
  f1,
  f2,
  f3;
assign
  g0 = \[0] ,
  h0 = \[1] ,
  i0 = \[2] ,
  k1 = ~o1 & (~n1 & (~m1 & ~l1)),
  k2 = ~o2 & (~n2 & (~m2 & ~l2)),
  l1 = (~f0 & p) | (f0 & ~p),
  l2 = (~\x  & h) | (\x  & ~h),
  m0 = ~k1 & ~c1,
  m1 = (~e0 & o) | (e0 & ~o),
  m2 = (~w & g) | (w & ~g),
  n1 = (~d0 & n) | (d0 & ~n),
  n2 = (~v & f) | (v & ~f),
  o0 = ~x1 & ~d1,
  o1 = (~c0 & m) | (c0 & ~m),
  o2 = (~u & e) | (u & ~e),
  p1 = f0 | ~p,
  p2 = \x  | ~h,
  \[0]  = ~\[1]  & ~\[2] ,
  q0 = ~k2 & ~e1,
  q1 = e0 | ~o,
  q2 = w | ~g,
  \[1]  = ~x0 & (~w0 & (~v0 & ~u0)),
  r1 = d0 | ~n,
  r2 = v | ~f,
  \[2]  = (~y0 & (~x0 & (~w0 & ~v0))) | ((~z0 & (~x0 & ~w0)) | ((~a1 & ~x0) | ~b1)),
  s0 = ~x2 & ~f1,
  s1 = c0 | ~m,
  s2 = u | ~e,
  u0 = (~m0 & c1) | (m0 & ~c1),
  v0 = (~o0 & d1) | (o0 & ~d1),
  w0 = (~q0 & e1) | (q0 & ~e1),
  x0 = (~s0 & f1) | (s0 & ~f1),
  x1 = ~b2 & (~a2 & (~z1 & ~y1)),
  x2 = ~b3 & (~a3 & (~z2 & ~y2)),
  y0 = m0 | ~c1,
  y1 = (~b0 & l) | (b0 & ~l),
  y2 = (~t & d) | (t & ~d),
  z0 = o0 | ~d1,
  z1 = (~a0 & k) | (a0 & ~k),
  z2 = (~s & c) | (s & ~c),
  a1 = q0 | ~e1,
  a2 = (~z & j) | (z & ~j),
  a3 = (~r & b) | (r & ~b),
  b1 = s0 | ~f1,
  b2 = (~y & i) | (y & ~i),
  b3 = (~q & a) | (q & ~a),
  c1 = (~p1 & (~o1 & (~n1 & ~m1))) | ((~q1 & (~o1 & ~n1)) | ((~r1 & ~o1) | ~s1)),
  c2 = b0 | ~l,
  c3 = t | ~d,
  d1 = (~c2 & (~b2 & (~a2 & ~z1))) | ((~d2 & (~b2 & ~a2)) | ((~e2 & ~b2) | ~f2)),
  d2 = a0 | ~k,
  d3 = s | ~c,
  e1 = (~p2 & (~o2 & (~n2 & ~m2))) | ((~q2 & (~o2 & ~n2)) | ((~r2 & ~o2) | ~s2)),
  e2 = z | ~j,
  e3 = r | ~b,
  f1 = (~c3 & (~b3 & (~a3 & ~z2))) | ((~d3 & (~b3 & ~a3)) | ((~e3 & ~b3) | ~f3)),
  f2 = y | ~i,
  f3 = q | ~a;
endmodule

