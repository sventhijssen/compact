// IWLS benchmark module "rot" printed on Wed May 29 16:09:27 2002
module rot(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, \x , y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2, b2, c2, d2, e2, f2, g2, h2, i2, j2, k2, l2, m2, n2, o2, p2, q2, r2, s2, t2, u2, v2, w2, x2, y2, z2, a3, b3, c3, d3, e3, f3, g3, h3, i3, j3, k3, l3, m3, n3, o3, p3, q3, r3, s3, t3, u3, v3, w3, x3, y3, z3, a4, b4, c4, d4, e4, f4, g4, h4, i4, j4, k4, l4, m4, n4, o4, p4, q4, r4, s4, t4, u4, v4, w4, x4, y4, z4, a5, b5, c5, d5, e5, f5, g5, h5, i5, j5, k5, l5, m5, n5, o5, p5, q5, r5, s5, t5, u5, v5, w5, x5, y5, z5, a6, b6, c6, d6, e6, f6, g6, h6, i6, j6, k6, l6, m6, n6, o6, p6, q6, r6, s6, t6, u6, v6, w6, x6, y6, z6, a7, b7, c7, d7, e7, f7, g7, h7, i7, j7, k7, l7, m7, n7, o7, p7, q7, r7, s7, t7, u7, v7, w7, x7, y7, z7, a8, b8, c8, d8, e8, f8, g8, h8);
input
  z0,
  z1,
  z2,
  z3,
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  t,
  u,
  v,
  w,
  \x ,
  y,
  z,
  a0,
  a1,
  a2,
  a3,
  a4,
  b0,
  b1,
  b2,
  b3,
  b4,
  c0,
  c1,
  c2,
  c3,
  c4,
  d0,
  d1,
  d2,
  d3,
  d4,
  e0,
  e1,
  e2,
  e3,
  e4,
  f0,
  f1,
  f2,
  f3,
  g0,
  g1,
  g2,
  g3,
  h0,
  h1,
  h2,
  h3,
  i0,
  i1,
  i2,
  i3,
  j0,
  j1,
  j2,
  j3,
  k0,
  k1,
  k2,
  k3,
  l0,
  l1,
  l2,
  l3,
  m0,
  m1,
  m2,
  m3,
  n0,
  n1,
  n2,
  n3,
  o0,
  o1,
  o2,
  o3,
  p0,
  p1,
  p2,
  p3,
  q0,
  q1,
  q2,
  q3,
  r0,
  r1,
  r2,
  r3,
  s0,
  s1,
  s2,
  s3,
  t0,
  t1,
  t2,
  t3,
  u0,
  u1,
  u2,
  u3,
  v0,
  v1,
  v2,
  v3,
  w0,
  w1,
  w2,
  w3,
  x0,
  x1,
  x2,
  x3,
  y0,
  y1,
  y2,
  y3;
output
  z4,
  z5,
  z6,
  z7,
  a5,
  a6,
  a7,
  a8,
  b5,
  b6,
  b7,
  b8,
  c5,
  c6,
  c7,
  c8,
  d5,
  d6,
  d7,
  d8,
  e5,
  e6,
  e7,
  e8,
  f4,
  f5,
  f6,
  f7,
  f8,
  g4,
  g5,
  g6,
  g7,
  g8,
  h4,
  h5,
  h6,
  h7,
  h8,
  i4,
  i5,
  i6,
  i7,
  j4,
  j5,
  j6,
  j7,
  k4,
  k5,
  k6,
  k7,
  l4,
  l5,
  l6,
  l7,
  m4,
  m5,
  m6,
  m7,
  n4,
  n5,
  n6,
  n7,
  o4,
  o5,
  o6,
  o7,
  p4,
  p5,
  p6,
  p7,
  q4,
  q5,
  q6,
  q7,
  r4,
  r5,
  r6,
  r7,
  s4,
  s5,
  s6,
  s7,
  t4,
  t5,
  t6,
  t7,
  u4,
  u5,
  u6,
  u7,
  v4,
  v5,
  v6,
  v7,
  w4,
  w5,
  w6,
  w7,
  x4,
  x5,
  x6,
  x7,
  y4,
  y5,
  y6,
  y7;
wire
  j13,
  j14,
  j15,
  j16,
  \[146] ,
  r12,
  \[148] ,
  r13,
  r14,
  r15,
  z12,
  z13,
  z14,
  z16,
  \[150] ,
  c13,
  c14,
  c15,
  c16,
  \[153] ,
  k13,
  k14,
  k15,
  k17,
  \[6] ,
  s12,
  \[158] ,
  s13,
  s14,
  s15,
  s16,
  \[159] ,
  \[161] ,
  d13,
  d14,
  d15,
  d16,
  d17,
  \[162] ,
  \[163] ,
  l12,
  l13,
  l14,
  l15,
  \[165] ,
  l17,
  t12,
  \[168] ,
  t13,
  t14,
  t15,
  \[171] ,
  e13,
  e14,
  e15,
  e16,
  \[174] ,
  m12,
  m13,
  m14,
  m15,
  m16,
  \[176] ,
  u12,
  u13,
  u14,
  u15,
  \[179] ,
  \[181] ,
  f13,
  f14,
  f15,
  f16,
  f17,
  \[182] ,
  \[183] ,
  \[200] ,
  \[107] ,
  \[201] ,
  n12,
  \[108] ,
  n13,
  n14,
  n15,
  \[185] ,
  \[202] ,
  \[109] ,
  v12,
  v13,
  v15,
  v16,
  \[110] ,
  \[112] ,
  \[113] ,
  \[190] ,
  \[114] ,
  g13,
  g14,
  g15,
  \[115] ,
  g16,
  \[117] ,
  o12,
  \[118] ,
  o13,
  o14,
  o15,
  o16,
  \[197] ,
  w12,
  w13,
  w15,
  w16,
  \[199] ,
  \[120] ,
  \[122] ,
  \[123] ,
  h13,
  h14,
  h15,
  \[125] ,
  h16,
  h17,
  \[126] ,
  \[127] ,
  p12,
  \[128] ,
  p13,
  p14,
  p15,
  p16,
  p17,
  \[129] ,
  x12,
  x13,
  x14,
  x15,
  \[130] ,
  \[131] ,
  a13,
  a14,
  a15,
  \[132] ,
  \[133] ,
  \[134] ,
  \[50] ,
  i13,
  i14,
  i15,
  \[135] ,
  i16,
  \[137] ,
  q12,
  q13,
  q14,
  q15,
  q16,
  y12,
  y13,
  y14,
  y15,
  y16,
  \[141] ,
  b13,
  b14,
  b15,
  b16;
assign
  z4 = c13,
  z5 = a14,
  z6 = x14,
  z7 = q15,
  j13 = l13 & k13,
  j14 = (\[131]  & (~g16 & r0)) | o16,
  j15 = h16 & ~s16,
  j16 = \[197]  & a2,
  \[146]  = \[123]  | (p | ~o),
  r12 = v16 & w1,
  \[148]  = ~b16 | n2,
  r13 = (~\[130]  & x13) | ((~p16 & j16) | ((~p16 & j0) | (p16 & i16))),
  r14 = (\[201]  & (~g16 & c3)) | (q14 & c3),
  r15 = (w16 & v16) | c4,
  z12 = (~y15 & (b & ~x15)) | ((y15 & (~b & ~x15)) | (x15 & d2)),
  z13 = (\[179]  & l3) | ~\[115] ,
  z14 = (y14 & (~y3 & (o1 & m1))) | ((y14 & (m1 & i1)) | ((e14 & (~y3 & o1)) | ((~y3 & (~l2 & o1)) | ((~y3 & (o1 & ~q)) | ((e14 & i1) | ((~l2 & i1) | (i1 & ~q))))))),
  z16 = (~v15 & (x14 & ~w0)) | ((v15 & (~x14 & ~z0)) | (z0 & w0)),
  \[150]  = z16 | p17,
  c13 = b4 & v0,
  c14 = (\[163]  & m2) | (m2 & m1),
  c15 = (~k1 & k17) | (~k17 & q3),
  c16 = (\[200]  & (\[126]  & ~g16)) | (\[126]  & (i3 & h3)),
  \[153]  = q16 | ~u2,
  k13 = (l2 & ~d1) | \[158] ,
  k14 = ~k2 & ~m0,
  k15 = (~\[197]  & ~h16) | s16,
  k17 = (~\[110]  & (~m2 & q)) | (\[182]  & \[110] ),
  \[6]  = ~o3,
  s12 = (\[134]  & (\[113]  & (\[107]  & (x15 & ~a)))) | ((\[134]  & (\[113]  & (\[107]  & (q16 & ~a)))) | ((\[113]  & (\[107]  & (x15 & (~o13 & ~h2)))) | ((\[113]  & (\[107]  & (x15 & (~o13 & ~f2)))) | ((\[113]  & (\[107]  & (q16 & (~o13 & ~h2)))) | ((\[113]  & (\[107]  & (q16 & (~o13 & ~f2)))) | ((~\[120]  & (\[107]  & (x15 & ~o13))) | (~\[120]  & (\[107]  & (q16 & ~o13))))))))),
  \[158]  = (l2 & p) | ((l2 & ~n) | ~\[123] ),
  s13 = p16 & (~i16 & ~o16),
  s14 = (\[201]  & d3) | (c3 & o0),
  s15 = ~w16 & (v16 & (x2 & ~w2)),
  s16 = (\[127]  & n1) | (\[122]  & n1),
  \[159]  = m2 & y1,
  \[161]  = ~y15 | ~b,
  d13 = (~d1 & c1) | (d1 & ~c1),
  d14 = \[181]  & w1,
  d15 = (~l1 & (k1 & k17)) | ((l1 & (~k1 & k17)) | (~k17 & r3)),
  d16 = (~i3 & h3) | ~\[141] ,
  d17 = ~\[130]  & ~\[126] ,
  \[162]  = ~d1 | ~c1,
  \[163]  = q2 | r0,
  l12 = (~\[183]  & j1) | (\[183]  & e0),
  l13 = (l2 & ~c1) | \[158] ,
  l14 = (~d16 & (m2 & ~k2)) | ((~i3 & (m2 & ~k2)) | ((p2 & ~k2) | k14)),
  l15 = (\[202]  & (\[125]  & (\[108]  & (~h16 & (a4 & l3))))) | ((\[202]  & (\[125]  & (\[114]  & (~h16 & a4)))) | ((\[125]  & (\[114]  & (~h16 & (p16 & a4)))) | ((\[125]  & (\[108]  & (~h16 & (i14 & a4)))) | ((\[202]  & (~q16 & (~u15 & a4))) | ((\[174]  & (\[125]  & (h16 & a4))) | ((s16 & (~q16 & (~u15 & a4))) | ((h16 & (~q16 & (~u15 & a4))) | ((p16 & (~q16 & (~u15 & a4))) | (\[125]  & (s16 & a4)))))))))),
  \[165]  = l3 | s,
  l17 = (\[181]  & (\[110]  & r0)) | (~\[110]  & (~m2 & p)),
  t12 = (~\[120]  & (~\[107]  & ~a)) | (t2 & a1),
  \[168]  = s16 | ~y3,
  t13 = (~\[150]  & j2) | (j16 & ~o3),
  t14 = (~\[150]  & j2) | (~\[146]  & ~k2),
  t15 = (~v16 & w2) | ~a4,
  \[171]  = \[109]  | ~c16,
  e13 = (~\[162]  & ~e1) | (\[162]  & e1),
  e14 = (~q2 & p2) | (q2 & ~p2),
  e15 = \[202]  & y3,
  e16 = (~d3 & (~c3 & ~b3)) | ((d3 & (l2 & o0)) | (~c3 & (l2 & o0))),
  \[174]  = \[133] ,
  m12 = (~y1 & p0) | (y1 & k1),
  m13 = ~\[162]  & (e1 & n),
  m14 = (y16 & h3) | (d17 | o16),
  m15 = \[176]  & ~s1,
  m16 = (~\[174]  & (~\[132]  & h16)) | ((~\[165]  & (~\[132]  & u2)) | ((~\[132]  & (~\[108]  & u2)) | ((~\[132]  & ~\[125] ) | ((v16 & u15) | (~w15 & ~x2))))),
  \[176]  = (w16 & v16) | (u15 | d4),
  u12 = (\[127]  & (~h2 & (~r1 & (~q1 & (~h1 & (~g1 & (~f1 & a))))))) | ((\[134]  & (\[127]  & (\[112]  & (~f17 & (~r1 & ~q1))))) | ((\[134]  & (\[127]  & (\[112]  & (~r1 & (~q1 & a))))) | ((\[134]  & (\[127]  & (~h2 & (~r1 & (~q1 & a))))) | ((~\[134]  & (\[112]  & (~h1 & (~g1 & ~f1)))) | (\[112]  & ~l2))))),
  u13 = (\[190]  & k0) | ((k0 & h0) | l2),
  u14 = \[179]  & ~p17,
  u15 = (~w16 & w2) | ((~v16 & x2) | (~x2 & w2)),
  \[179]  = t0 & g0,
  \[181]  = m2 & (~y1 & x1),
  f13 = j13 & h13,
  f14 = (\[163]  & m2) | (p2 & m2),
  f15 = ~u15 & ~m1,
  f16 = (\[200]  & \[129] ) | ((\[129]  & f3) | (\[129]  & e3)),
  f17 = (~h2 & (~g2 & f2)) | (h2 & (~g2 & ~f2)),
  \[182]  = \[159]  & ~x1,
  \[183]  = y | ~\x ,
  \[200]  = d16 & m3,
  \[107]  = ~t2 | t1,
  \[201]  = ~o0,
  n12 = u15 | v2,
  \[108]  = (b2 & ~s1) | ~s0,
  n13 = (\[199]  & ~\[127] ) | (\[199]  & b1),
  n14 = (~y16 & (~i3 & h3)) | ((y16 & i3) | d17),
  n15 = \[176]  & ~\[127] ,
  \[185]  = ~y | \x ,
  \[202]  = e4 & i1,
  \[109]  = (~s0 & h0) | (s0 & u),
  v12 = (h17 & (p12 & ~a)) | (f0 & ~a),
  v13 = (~\[153]  & l0) | ((~j16 & l0) | ((~s0 & l0) | \[113] )),
  v15 = ~x0 & ~w0,
  v16 = \[159]  & x1,
  \[110]  = ~q2 | ~p2,
  \[112]  = (h2 & (~q & (~p & ~o))) | o0,
  \[113]  = (f17 & l2) | z1,
  \[190]  = \[118]  | ~j16,
  \[114]  = (\[108]  & s) | ~u2,
  g13 = k13 & i13,
  g14 = (~p0 & l17) | (~l17 & v3),
  g15 = \[182]  | i1,
  \[115]  = ~\[150]  | ~j2,
  g16 = h17 & r1,
  \[117]  = ~f0 | ~a,
  o12 = (~s0 & (u2 & (h0 & ~g0))) | ((s0 & (u2 & (u & ~t))) | u15),
  \[118]  = a3 | z2,
  o13 = (~q13 & (~p13 & ~l2)) | a,
  o14 = (~d16 & z2) | ((~c16 & z2) | ~\[171] ),
  o15 = (~p3 & r) | ((k3 & r) | (s2 & u0)),
  o16 = ~l3 & (t0 & (h0 & ~g0)),
  \[197]  = t3 | (o3 | n3),
  w12 = (x15 & (~o12 & (~s0 & i0))) | ((x15 & (~o12 & (s0 & v))) | ((~b16 & (~x15 & n2)) | ((~\[148]  & ~x15) | ((\[137]  & x15) | (~\[133]  & x15))))),
  w13 = (\[141]  & (~\[123]  & (~o16 & (p & ~o)))) | ((~\[123]  & (~o16 & (p2 & p))) | ((\[181]  & (~o16 & ~w1)) | (~o16 & m0))),
  w15 = (~w2 & u15) | (~w2 & ~x2),
  w16 = (~\[109]  & (x2 & (~w2 & (u2 & (~d0 & ~m))))) | ((~\[109]  & (x2 & (~w2 & (u2 & (d0 & ~k))))) | ((~\[109]  & (u3 & (u2 & ~h))) | ((u3 & ~i) | ((~d0 & ~l) | ((d0 & ~j) | ~g))))),
  \[199]  = ~f | (~e | ~d),
  \[120]  = h2 | f2,
  \[122]  = u15 | ~b2,
  \[123]  = ~l2 | q,
  h13 = l13 & i13,
  h14 = (~q0 & (p0 & l17)) | ((q0 & (~p0 & l17)) | (~l17 & w3)),
  h15 = (x15 & u2) | ((~l3 & s) | h16),
  \[125]  = (~\[168]  & ~u15) | ~n12,
  h16 = ~g16 & (f16 & g3),
  h17 = (\[120]  & (\[113]  & (o2 & (~s1 & (r1 & ~p1))))) | (~\[127]  & (\[120]  & (\[113]  & (o2 & ~p1)))),
  \[126]  = \[118]  | e16,
  \[127]  = ~s1 | r1,
  p12 = (\[109]  & u2) | (u15 & c2),
  \[128]  = ~h17 | p12,
  p13 = (~q13 & (~l2 & ~g2)) | (~q13 & f2),
  p14 = (~\[171]  & (~s0 & i0)) | ((~\[171]  & (s0 & v)) | ((\[171]  & (~g16 & a3)) | ((\[171]  & (o14 & a3)) | (d16 & c16)))),
  p15 = p3 & j3,
  p16 = (\[135]  & (\[115]  & (j16 & (m0 & (l0 & k0))))) | (\[115]  & (m0 & (l0 & (k0 & j0)))),
  p17 = (~z16 & (~v15 & (u1 & (y0 & ~x0)))) | ((~z16 & (~x14 & (u1 & (~y0 & x0)))) | ((z16 & (u1 & (y0 & x0))) | (v15 & (x14 & u1)))),
  \[129]  = \[122]  | ~v1,
  x12 = (\[200]  & (~\[133]  & (x15 & (~i3 & f3)))) | ((\[200]  & (~\[133]  & (x15 & (i3 & e3)))) | ((~\[133]  & (x15 & (f3 & e3))) | ((\[148]  & (~x15 & o2)) | (\[137]  & x15)))),
  x13 = p16 & n3,
  x14 = ~z0 & ~y0,
  x15 = ~q16 & m16,
  a5 = m2,
  a6 = b14,
  a7 = y0,
  a8 = r15,
  b5 = d13,
  b6 = c14,
  b7 = z0,
  b8 = s15,
  c5 = e13,
  c6 = d14,
  c7 = y14,
  c8 = t15,
  d5 = f13,
  d6 = \[50] ,
  d7 = z14,
  d8 = u15,
  e5 = g13,
  e6 = e14,
  e7 = a15,
  e8 = v15,
  \[130]  = ~t0 | h0,
  f4 = l12,
  f5 = h13,
  f6 = f14,
  f7 = b15,
  f8 = w0,
  \[131]  = \[110]  | ~l2,
  g4 = m12,
  g5 = i13,
  g6 = g14,
  g7 = c15,
  a13 = (~\[161]  & (~x15 & ~c)) | ((\[161]  & (~x15 & c)) | (x15 & e2)),
  g8 = x0,
  a14 = ~\[135]  | (u15 | (k2 | i2)),
  a15 = \[165]  & (e15 & z3),
  \[132]  = u15 | z3,
  h4 = n12,
  h5 = j13,
  h6 = h14,
  h7 = d15,
  h8 = w15,
  \[133]  = ~f16 | ~y2,
  i4 = o12,
  i5 = k13,
  i6 = i14,
  i7 = e15,
  \[134]  = ~l2 | ~g2,
  \[50]  = ~p2,
  j4 = p12,
  j5 = l13,
  j6 = j14,
  j7 = f15,
  i13 = (l2 & ~e1) | \[158] ,
  i14 = p16 & l3,
  i15 = ~h16 & ~k15,
  \[135]  = \[130]  | ~n3,
  i16 = (\[179]  & (p17 & (j16 & ~l2))) | ((\[153]  & (j16 & (~l3 & t0))) | ((~\[190]  & (~\[130]  & ~l3)) | ((\[132]  & ~\[109] ) | (d16 & ~y16)))),
  k4 = s3,
  k5 = l2,
  k6 = k14,
  k7 = g15,
  l4 = \[6] ,
  l5 = m13,
  l6 = l14,
  l7 = h15,
  \[137]  = (~o12 & n12) | (o12 & ~n12),
  m4 = t3,
  m5 = n13,
  m6 = m14,
  m7 = i15,
  q12 = (\[181]  & (\[110]  & r0)) | ((\[182]  & m13) | ((\[182]  & ~n) | (v16 & ~r12))),
  q13 = (~l2 & ~h2) | ((l2 & f2) | ~\[134] ),
  q14 = \[201]  & b3,
  q15 = (~d0 & k) | (d0 & m),
  q16 = \[128]  & (\[117]  & r2),
  n4 = q12,
  n5 = o13,
  n6 = n14,
  n7 = j15,
  o4 = r12,
  o5 = p13,
  o6 = o14,
  o7 = k15,
  p4 = s12,
  p5 = q13,
  p6 = p14,
  p7 = l15,
  y12 = (\[128]  & (\[117]  & (~y15 & m16))) | ((\[128]  & (\[117]  & (b16 & m16))) | ((~y15 & q16) | (b16 & q16))),
  y13 = (\[179]  & (p17 & ~l2)) | (\[146]  & k2),
  y14 = (\[131]  & (~h17 & (~y3 & o1))) | ((\[131]  & (~y3 & (~s1 & o1))) | ((~h17 & (~y3 & (o1 & ~q))) | ((~y3 & (~s1 & (o1 & ~q))) | ((\[131]  & (~h17 & m1)) | ((\[131]  & (~s1 & m1)) | ((~h17 & (m1 & ~q)) | (~s1 & (m1 & ~q)))))))),
  y15 = (~\[199]  & a) | ((\[127]  & a) | (~n & a)),
  y16 = (~\[126]  & (~g16 & m3)) | (~\[126]  & (i3 & h3)),
  q4 = t12,
  q5 = r13,
  q6 = q14,
  q7 = m15,
  r4 = u12,
  r5 = s13,
  r6 = r14,
  r7 = n15,
  s4 = v12,
  s5 = t13,
  s6 = s14,
  s7 = w,
  t4 = w12,
  t5 = u13,
  t6 = t14,
  t7 = z,
  u4 = x12,
  u5 = v13,
  u6 = u14,
  u7 = a0,
  v4 = y12,
  v5 = w13,
  v6 = x14,
  v7 = b0,
  \[141]  = ~i3 | h3,
  w4 = z12,
  w5 = x13,
  w6 = y0,
  w7 = c0,
  b13 = (~x3 & v0) | a,
  b14 = (~\[185]  & e0) | (\[185]  & n0),
  b15 = (q2 & m2) | ((p2 & m2) | (m2 & m1)),
  b16 = (o2 & y15) | (n2 & y15),
  x4 = a13,
  x5 = y13,
  x6 = v15,
  x7 = o15,
  y4 = b13,
  y5 = z13,
  y6 = w0,
  y7 = p15;
endmodule

