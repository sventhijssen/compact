module s349(VDD,CK,A0,A1,A2,A3,B0,B1,B2,B3,CNTVCO2,CNTVCON2,P0,P1,P2,P3,P4,
  P5,P6,P7,READY,START);
input VDD,CK,START,B0,B1,B2,B3,A0,A1,A2,A3;
output CNTVCO2,CNTVCON2,READY,P0,P1,P2,P3,P4,P5,P6,P7;

  wire CT2,CNTVG3VD,CT1,CNTVG2VD,CT0,CNTVG1VD,ACVQN3,ACVG4VD1,ACVQN2,ACVG3VD1,
    ACVQN1,ACVG2VD1,ACVQN0,ACVG1VD1,MRVQN3,MRVG4VD,MRVQN2,MRVG3VD,MRVQN1,
    MRVG2VD,MRVQN0,MRVG1VD,AX3,AM3,AX2,AM2,AX1,AM1,AX0,AM0,READYN,CT1N,
    CNTVG3VQN,CNTVG2VQN,CNTVCO0,CNTVG1VQN,CNTVCON0,CNTVG1VD1,S3,ADDVG4VSN,CO,
    ADDVG4VCN,S2,ADDVG3VSN,ADDVC3,ADDVG3VCN,S1,ADDVG2VSN,ADDVC2,ADDVG2VCN,
    ADDVC1,ADDVG1VCN,S0,ADDVG1VP,AD0,AD0N,AD1,AD1N,AD2,AD2N,AD3,AD3N,ACVPCN,
    SMVG5VS0P,SMVS0N,SM3,SMVG5VX,SMVG4VS0P,SM2,SMVG4VX,SMVG3VS0P,SM1,SMVG3VX,
    SMVG2VS0P,SM0,SMVG2VX,ADSH,MRVSHLDN,BMVG5VS0P,BMVS0N,BM3,BMVG5VX,BMVG4VS0P,
    BM2,BMVG4VX,BMVG3VS0P,BM1,BMVG3VX,BMVG2VS0P,BM0,BMVG2VX,AMVG5VS0P,AMVS0N,
    AMVG5VX,AMVG4VS0P,AMVG4VX,AMVG3VS0P,AMVG3VX,AMVG2VS0P,AMVG2VX,IINIIT,
    ADDVG4VCNVAD4NF,ADDVG4VCNVAD3NF,ADDVG4VCNVOR2NF,ADDVG4VCNVAD2NF,
    ADDVG4VCNVOR1NF,ADDVG4VCNVAD1NF,ADDVG3VCNVAD4NF,ADDVG3VCNVAD3NF,
    ADDVG3VCNVOR2NF,ADDVG3VCNVAD2NF,ADDVG3VCNVOR1NF,ADDVG3VCNVAD1NF,
    ADDVG2VCNVAD4NF,ADDVG2VCNVAD3NF,ADDVG2VCNVOR2NF,ADDVG2VCNVAD2NF,
    ADDVG2VCNVOR1NF,ADDVG2VCNVAD1NF,SMVG5VG1VAD2NF,SMVG5VG1VAD1NF,
    SMVG4VG1VAD2NF,SMVG4VG1VAD1NF,SMVG3VG1VAD2NF,SMVG3VG1VAD1NF,SMVG2VG1VAD2NF,
    SMVG2VG1VAD1NF,MRVG4VDVAD2NF,MRVG4VDVAD1NF,MRVG3VDVAD2NF,MRVG3VDVAD1NF,
    MRVG2VDVAD2NF,MRVG2VDVAD1NF,MRVG1VDVAD2NF,MRVG1VDVAD1NF,BMVG5VG1VAD2NF,
    BMVG5VG1VAD1NF,BMVG4VG1VAD2NF,BMVG4VG1VAD1NF,BMVG3VG1VAD2NF,BMVG3VG1VAD1NF,
    BMVG2VG1VAD2NF,BMVG2VG1VAD1NF,AMVG5VG1VAD2NF,AMVG5VG1VAD1NF,AMVG4VG1VAD2NF,
    AMVG4VG1VAD1NF,AMVG3VG1VAD2NF,AMVG3VG1VAD1NF,AMVG2VG1VAD2NF,AMVG2VG1VAD1NF,
    CNTVG3VG2VOR1NF,CNTVG3VD1,CNTVG2VG2VOR1NF,CNTVG2VD1,CNTVG1VG2VOR1NF,
    ADDVG1VPVOR1NF,CNTVCO1,CNTVG3VZ,CNTVG3VZ1,CNTVCON1,CNTVG2VZ,CNTVG2VZ1,
    CNTVG1VZ,CNTVG1VZ1;

  FD1 DFF_0(CK,CT2,CNTVG3VD);
  FD1 DFF_1(CK,CT1,CNTVG2VD);
  FD1 DFF_2(CK,CT0,CNTVG1VD);
  FD1 DFF_3(CK,ACVQN3,ACVG4VD1);
  FD1 DFF_4(CK,ACVQN2,ACVG3VD1);
  FD1 DFF_5(CK,ACVQN1,ACVG2VD1);
  FD1 DFF_6(CK,ACVQN0,ACVG1VD1);
  FD1 DFF_7(CK,MRVQN3,MRVG4VD);
  FD1 DFF_8(CK,MRVQN2,MRVG3VD);
  FD1 DFF_9(CK,MRVQN1,MRVG2VD);
  FD1 DFF_10(CK,MRVQN0,MRVG1VD);
  FD1 DFF_11(CK,AX3,AM3);
  FD1 DFF_12(CK,AX2,AM2);
  FD1 DFF_13(CK,AX1,AM1);
  FD1 DFF_14(CK,AX0,AM0);
  IV  NOT_0(READY,READYN);
  IV  NOT_1(CT1N,CT1);
  IV  NOT_2(CNTVG3VQN,CT2);
  IV  NOT_3(CNTVG2VQN,CT1);
  IV  NOT_4(CNTVCO0,CNTVG1VQN);
  IV  NOT_5(CNTVCON0,CT0);
  IV  NOT_6(CNTVG1VQN,CT0);
  IV  NOT_7(CNTVG1VD1,READY);
  IV  NOT_8(S3,ADDVG4VSN);
  IV  NOT_9(CO,ADDVG4VCN);
  IV  NOT_10(S2,ADDVG3VSN);
  IV  NOT_11(ADDVC3,ADDVG3VCN);
  IV  NOT_12(S1,ADDVG2VSN);
  IV  NOT_13(ADDVC2,ADDVG2VCN);
  IV  NOT_14(ADDVC1,ADDVG1VCN);
  IV  NOT_15(S0,ADDVG1VP);
  IV  NOT_16(AD0,AD0N);
  IV  NOT_17(AD1,AD1N);
  IV  NOT_18(AD2,AD2N);
  IV  NOT_19(AD3,AD3N);
  IV  NOT_20(ACVPCN,START);
  IV  NOT_21(P7,ACVQN3);
  IV  NOT_22(P6,ACVQN2);
  IV  NOT_23(P5,ACVQN1);
  IV  NOT_24(P4,ACVQN0);
  IV  NOT_25(SMVG5VS0P,SMVS0N);
  IV  NOT_26(SM3,SMVG5VX);
  IV  NOT_27(SMVG4VS0P,SMVS0N);
  IV  NOT_28(SM2,SMVG4VX);
  IV  NOT_29(SMVG3VS0P,SMVS0N);
  IV  NOT_30(SM1,SMVG3VX);
  IV  NOT_31(SMVG2VS0P,SMVS0N);
  IV  NOT_32(SM0,SMVG2VX);
  IV  NOT_33(SMVS0N,ADSH);
  IV  NOT_34(MRVSHLDN,ADSH);
  IV  NOT_35(P3,MRVQN3);
  IV  NOT_36(P2,MRVQN2);
  IV  NOT_37(P1,MRVQN1);
  IV  NOT_38(P0,MRVQN0);
  IV  NOT_39(BMVG5VS0P,BMVS0N);
  IV  NOT_40(BM3,BMVG5VX);
  IV  NOT_41(BMVG4VS0P,BMVS0N);
  IV  NOT_42(BM2,BMVG4VX);
  IV  NOT_43(BMVG3VS0P,BMVS0N);
  IV  NOT_44(BM1,BMVG3VX);
  IV  NOT_45(BMVG2VS0P,BMVS0N);
  IV  NOT_46(BM0,BMVG2VX);
  IV  NOT_47(BMVS0N,READYN);
  IV  NOT_48(AMVG5VS0P,AMVS0N);
  IV  NOT_49(AM3,AMVG5VX);
  IV  NOT_50(AMVG4VS0P,AMVS0N);
  IV  NOT_51(AM2,AMVG4VX);
  IV  NOT_52(AMVG3VS0P,AMVS0N);
  IV  NOT_53(AM1,AMVG3VX);
  IV  NOT_54(AMVG2VS0P,AMVS0N);
  IV  NOT_55(AM0,AMVG2VX);
  IV  NOT_56(AMVS0N,IINIIT);
  AN3 AND3_0(ADDVG4VCNVAD4NF,ADDVC3,AD3,P7);
  AN2 AND2_0(ADDVG4VCNVAD3NF,ADDVG4VCNVOR2NF,ADDVG4VCN);
  AN2 AND2_1(ADDVG4VCNVAD2NF,ADDVC3,ADDVG4VCNVOR1NF);
  AN2 AND2_2(ADDVG4VCNVAD1NF,AD3,P7);
  AN3 AND3_1(ADDVG3VCNVAD4NF,ADDVC2,AD2,P6);
  AN2 AND2_3(ADDVG3VCNVAD3NF,ADDVG3VCNVOR2NF,ADDVG3VCN);
  AN2 AND2_4(ADDVG3VCNVAD2NF,ADDVC2,ADDVG3VCNVOR1NF);
  AN2 AND2_5(ADDVG3VCNVAD1NF,AD2,P6);
  AN3 AND3_2(ADDVG2VCNVAD4NF,ADDVC1,AD1,P5);
  AN2 AND2_6(ADDVG2VCNVAD3NF,ADDVG2VCNVOR2NF,ADDVG2VCN);
  AN2 AND2_7(ADDVG2VCNVAD2NF,ADDVC1,ADDVG2VCNVOR1NF);
  AN2 AND2_8(ADDVG2VCNVAD1NF,AD1,P5);
  AN2 AND2_9(SMVG5VG1VAD2NF,SMVG5VS0P,CO);
  AN2 AND2_10(SMVG5VG1VAD1NF,SMVS0N,P7);
  AN2 AND2_11(SMVG4VG1VAD2NF,SMVG4VS0P,S3);
  AN2 AND2_12(SMVG4VG1VAD1NF,SMVS0N,P6);
  AN2 AND2_13(SMVG3VG1VAD2NF,SMVG3VS0P,S2);
  AN2 AND2_14(SMVG3VG1VAD1NF,SMVS0N,P5);
  AN2 AND2_15(SMVG2VG1VAD2NF,SMVG2VS0P,S1);
  AN2 AND2_16(SMVG2VG1VAD1NF,SMVS0N,P4);
  AN2 AND2_17(MRVG4VDVAD2NF,MRVSHLDN,BM3);
  AN2 AND2_18(MRVG4VDVAD1NF,ADSH,S0);
  AN2 AND2_19(MRVG3VDVAD2NF,MRVSHLDN,BM2);
  AN2 AND2_20(MRVG3VDVAD1NF,ADSH,P3);
  AN2 AND2_21(MRVG2VDVAD2NF,MRVSHLDN,BM1);
  AN2 AND2_22(MRVG2VDVAD1NF,ADSH,P2);
  AN2 AND2_23(MRVG1VDVAD2NF,MRVSHLDN,BM0);
  AN2 AND2_24(MRVG1VDVAD1NF,ADSH,P1);
  AN2 AND2_25(BMVG5VG1VAD2NF,BMVG5VS0P,B3);
  AN2 AND2_26(BMVG5VG1VAD1NF,BMVS0N,P3);
  AN2 AND2_27(BMVG4VG1VAD2NF,BMVG4VS0P,B2);
  AN2 AND2_28(BMVG4VG1VAD1NF,BMVS0N,P2);
  AN2 AND2_29(BMVG3VG1VAD2NF,BMVG3VS0P,B1);
  AN2 AND2_30(BMVG3VG1VAD1NF,BMVS0N,P1);
  AN2 AND2_31(BMVG2VG1VAD2NF,BMVG2VS0P,B0);
  AN2 AND2_32(BMVG2VG1VAD1NF,BMVS0N,P0);
  AN2 AND2_33(AMVG5VG1VAD2NF,AMVG5VS0P,A3);
  AN2 AND2_34(AMVG5VG1VAD1NF,AMVS0N,AX3);
  AN2 AND2_35(AMVG4VG1VAD2NF,AMVG4VS0P,A2);
  AN2 AND2_36(AMVG4VG1VAD1NF,AMVS0N,AX2);
  AN2 AND2_37(AMVG3VG1VAD2NF,AMVG3VS0P,A1);
  AN2 AND2_38(AMVG3VG1VAD1NF,AMVS0N,AX1);
  AN2 AND2_39(AMVG2VG1VAD2NF,AMVG2VS0P,A0);
  AN2 AND2_40(AMVG2VG1VAD1NF,AMVS0N,AX0);
  OR2 OR2_0(CNTVG3VG2VOR1NF,CT2,CNTVG3VD1);
  OR2 OR2_1(CNTVG2VG2VOR1NF,CT1,CNTVG2VD1);
  OR2 OR2_2(CNTVG1VG2VOR1NF,CT0,CNTVG1VD1);
  OR3 OR3_0(ADDVG4VCNVOR2NF,ADDVC3,AD3,P7);
  OR2 OR2_3(ADDVG4VCNVOR1NF,AD3,P7);
  OR3 OR3_1(ADDVG3VCNVOR2NF,ADDVC2,AD2,P6);
  OR2 OR2_4(ADDVG3VCNVOR1NF,AD2,P6);
  OR3 OR3_2(ADDVG2VCNVOR2NF,ADDVC1,AD1,P5);
  OR2 OR2_5(ADDVG2VCNVOR1NF,AD1,P5);
  OR2 OR2_6(ADDVG1VPVOR1NF,AD0,P4);
  ND3 NAND3_0(READYN,CT0,CT1N,CT2);
  ND2 NAND2_0(CNTVCON2,CT2,CNTVCO1);
  ND2 NAND2_1(CNTVG3VZ,CNTVG3VG2VOR1NF,CNTVG3VZ1);
  ND2 NAND2_2(CNTVG3VZ1,CT2,CNTVG3VD1);
  ND2 NAND2_3(CNTVCON1,CT1,CNTVCO0);
  ND2 NAND2_4(CNTVG2VZ,CNTVG2VG2VOR1NF,CNTVG2VZ1);
  ND2 NAND2_5(CNTVG2VZ1,CT1,CNTVG2VD1);
  ND2 NAND2_6(CNTVG1VZ,CNTVG1VG2VOR1NF,CNTVG1VZ1);
  ND2 NAND2_7(CNTVG1VZ1,CT0,CNTVG1VD1);
  ND2 NAND2_8(ADDVG1VP,ADDVG1VPVOR1NF,ADDVG1VCN);
  ND2 NAND2_9(ADDVG1VCN,AD0,P4);
  ND2 NAND2_10(AD0N,P0,AX0);
  ND2 NAND2_11(AD1N,P0,AX1);
  ND2 NAND2_12(AD2N,P0,AX2);
  ND2 NAND2_13(AD3N,P0,AX3);
  ND2 NAND2_14(ACVG4VD1,ACVPCN,SM3);
  ND2 NAND2_15(ACVG3VD1,ACVPCN,SM2);
  ND2 NAND2_16(ACVG2VD1,ACVPCN,SM1);
  ND2 NAND2_17(ACVG1VD1,ACVPCN,SM0);
  NR2 NOR2_0(ADSH,READY,IINIIT);
  NR3 NOR3_0(IINIIT,CT0,CT1,CT2);
  NR2 NOR2_1(CNTVCO2,CNTVG3VQN,CNTVCON1);
  NR2 NOR2_2(CNTVG3VD,CNTVG3VZ,START);
  NR2 NOR2_3(CNTVG3VD1,READY,CNTVCON1);
  NR2 NOR2_4(CNTVCO1,CNTVG2VQN,CNTVCON0);
  NR2 NOR2_5(CNTVG2VD,CNTVG2VZ,START);
  NR2 NOR2_6(CNTVG2VD1,READY,CNTVCON0);
  NR2 NOR2_7(CNTVG1VD,CNTVG1VZ,START);
  NR2 NOR2_8(ADDVG4VSN,ADDVG4VCNVAD4NF,ADDVG4VCNVAD3NF);
  NR2 NOR2_9(ADDVG4VCN,ADDVG4VCNVAD2NF,ADDVG4VCNVAD1NF);
  NR2 NOR2_10(ADDVG3VSN,ADDVG3VCNVAD4NF,ADDVG3VCNVAD3NF);
  NR2 NOR2_11(ADDVG3VCN,ADDVG3VCNVAD2NF,ADDVG3VCNVAD1NF);
  NR2 NOR2_12(ADDVG2VSN,ADDVG2VCNVAD4NF,ADDVG2VCNVAD3NF);
  NR2 NOR2_13(ADDVG2VCN,ADDVG2VCNVAD2NF,ADDVG2VCNVAD1NF);
  NR2 NOR2_14(SMVG5VX,SMVG5VG1VAD2NF,SMVG5VG1VAD1NF);
  NR2 NOR2_15(SMVG4VX,SMVG4VG1VAD2NF,SMVG4VG1VAD1NF);
  NR2 NOR2_16(SMVG3VX,SMVG3VG1VAD2NF,SMVG3VG1VAD1NF);
  NR2 NOR2_17(SMVG2VX,SMVG2VG1VAD2NF,SMVG2VG1VAD1NF);
  NR2 NOR2_18(MRVG4VD,MRVG4VDVAD2NF,MRVG4VDVAD1NF);
  NR2 NOR2_19(MRVG3VD,MRVG3VDVAD2NF,MRVG3VDVAD1NF);
  NR2 NOR2_20(MRVG2VD,MRVG2VDVAD2NF,MRVG2VDVAD1NF);
  NR2 NOR2_21(MRVG1VD,MRVG1VDVAD2NF,MRVG1VDVAD1NF);
  NR2 NOR2_22(BMVG5VX,BMVG5VG1VAD2NF,BMVG5VG1VAD1NF);
  NR2 NOR2_23(BMVG4VX,BMVG4VG1VAD2NF,BMVG4VG1VAD1NF);
  NR2 NOR2_24(BMVG3VX,BMVG3VG1VAD2NF,BMVG3VG1VAD1NF);
  NR2 NOR2_25(BMVG2VX,BMVG2VG1VAD2NF,BMVG2VG1VAD1NF);
  NR2 NOR2_26(AMVG5VX,AMVG5VG1VAD2NF,AMVG5VG1VAD1NF);
  NR2 NOR2_27(AMVG4VX,AMVG4VG1VAD2NF,AMVG4VG1VAD1NF);
  NR2 NOR2_28(AMVG3VX,AMVG3VG1VAD2NF,AMVG3VG1VAD1NF);
  NR2 NOR2_29(AMVG2VX,AMVG2VG1VAD2NF,AMVG2VG1VAD1NF);

endmodule
