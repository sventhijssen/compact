module foobar(y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0);
input a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0;
output y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1;
not(y0, q10);
not(z0, n10);
not(t_0, c31);
not(t_1, d23);
or(a1, t_0, t_1);
not(t_2, f44);
not(t_3, e44);
or(b1, t_2, t_3);
not(t_4, n47);
not(t_5, o47);
or(c1, t_4, t_5);
and(d1, w46, f47);
not(e1, g50);
or(f1, x52, z53);
and(g1, t55, s56);
and(h1, t56, l57);
and(i1, t58, n59);
and(j1, p60, w60);
and(k1, h61, t61);
and(l1, b61, m61);
and(m1, z60, k61);
and(p1, q61, e62);
not(q1, d63);
not(r1, t63);
and(s1, t65, u65);
not(t_6, w65);
not(t_7, v65);
or(t1, t_6, t_7);
buf(o2, v0);
buf(p2, u0);
buf(q2, k0);
buf(r2, j0);
or(s2, j0, i0);
buf(t2, i0);
buf(u2, h0);
buf(v2, g0);
buf(w2, f0);
buf(x2, e0);
buf(y2, d0);
not(z2, a0);
not(a3, z);
buf(b3, y);
buf(c3, x);
not(d3, n);
buf(e3, n);
buf(f3, m);
not(g3, m);
not(h3, m);
buf(i3, m);
buf(j3, l);
buf(k3, l);
not(l3, l);
buf(m3, l);
not(n3, l);
buf(o3, l);
not(p3, k);
buf(q3, k);
not(r3, k);
buf(s3, k);
buf(t3, j);
not(u3, j);
buf(v3, j);
buf(w3, i);
not(x3, i);
buf(y3, i);
buf(z3, i);
not(a4, i);
buf(b4, i);
buf(c4, h);
buf(d4, h);
not(e4, h);
buf(f4, h);
not(g4, h);
buf(h4, h);
not(i4, g);
buf(j4, g);
not(k4, g);
buf(l4, g);
not(m4, f);
buf(n4, f);
or(o4, f, e);
not(p4, e);
not(q4, d);
or(r4, d, w0);
not(s4, d);
buf(t4, d);
not(u4, d);
and(v4, d, e);
not(w4, c);
not(x4, c);
and(y4, c, x);
not(t_8, z);
not(t_9, c);
or(z4, t_8, t_9);
and(a5, c, z);
not(b5, c);
not(c5, c);
not(d5, c);
buf(e5, c);
not(f5, b);
buf(g5, b);
and(h5, b, c);
not(t_10, d);
not(t_11, c);
not(t_12, a);
or(i5, t_10, t_11, t_12);
not(t_13, b);
not(t_14, a);
or(j5, t_13, t_14);
not(k5, a);
buf(l5, a);
not(m5, a);
buf(n5, a);
or(o5, o2, z2);
not(t_15, z2);
not(t_16, o2);
and(p5, t_15, t_16);
not(q5, p2);
not(r5, q2);
not(t_17, e3);
not(t_18, k0);
or(s5, t_17, t_18);
not(t5, r2);
not(t_19, i3);
not(t_20, j0);
or(u5, t_19, t_20);
not(v5, t2);
not(t_21, o3);
not(t_22, i0);
or(w5, t_21, t_22);
and(x5, h0, s2);
not(y5, u2);
not(t_23, s3);
not(t_24, h0);
or(z5, t_23, t_24);
not(a6, v2);
not(t_25, t3);
not(t_26, g0);
or(b6, t_25, t_26);
not(c6, w2);
not(t_27, z3);
not(t_28, f0);
or(d6, t_27, t_28);
not(e6, x2);
not(t_29, h4);
not(t_30, e0);
or(f6, t_29, t_30);
not(g6, y2);
not(t_31, l4);
not(t_32, d0);
or(h6, t_31, t_32);
or(i6, b3, b5);
not(t_33, b5);
not(t_34, b3);
and(j6, t_33, t_34);
not(k6, c3);
or(l6, w, x4);
buf(m6, d3);
buf(n6, f3);
buf(o6, f3);
and(p6, p3, l3, g3);
not(t_35, g3);
not(t_36, l3);
not(t_37, p3);
or(q6, t_35, t_36, t_37);
buf(r6, h3);
not(t_38, h3);
not(t_39, n3);
or(s6, t_38, t_39);
not(t6, j3);
not(u6, k3);
buf(v6, n3);
buf(w6, r3);
buf(x6, u3);
not(t_40, v3);
not(t_41, b4);
or(y6, t_40, t_41);
buf(z6, w3);
buf(a7, w3);
and(b7, i4, e4, x3);
not(t_42, x3);
not(t_43, e4);
not(t_44, i4);
or(c7, t_42, t_43, t_44);
buf(d7, a4);
not(t_45, a4);
not(t_46, g4);
or(e7, t_45, t_46);
not(f7, c4);
not(g7, d4);
buf(h7, g4);
not(i7, j4);
buf(j7, k4);
not(t_47, f);
not(t_48, d5);
not(t_49, g5);
or(k7, t_47, t_48, t_49);
buf(l7, m4);
buf(m7, m4);
and(n7, k5, n4, p4);
and(o7, m5, n4);
and(p7, k5, o4);
buf(q7, p4);
not(r7, r4);
not(s7, r4);
not(t7, r4);
not(u7, r4);
not(v7, r4);
not(w7, r4);
not(x7, r4);
not(y7, r4);
buf(z7, s4);
buf(a8, s4);
buf(b8, t4);
not(c8, v4);
not(d8, v4);
buf(e8, y4);
not(f8, y4);
or(g8, c, u4);
not(h8, c5);
not(i8, c5);
not(j8, c5);
not(k8, c5);
not(l8, c5);
not(m8, c5);
not(n8, c5);
not(o8, c5);
and(p8, m5, g5, d5);
and(q8, n5, f5, e5);
not(t_50, e5);
not(t_51, f5);
not(t_52, n5);
or(r8, t_50, t_51, t_52);
not(t_53, f5);
not(t_54, n5);
or(s8, t_53, t_54);
buf(t8, g5);
not(u8, h5);
or(v8, a, q4);
or(w8, a, w4);
and(x8, j5, i5);
buf(y8, l5);
buf(z8, p5);
not(t_55, t5);
not(t_56, q2);
or(a9, t_55, t_56);
and(b9, z5, w5, u5, s5);
not(t_57, r5);
not(t_58, r2);
or(c9, t_57, t_58);
and(d9, i0, y7);
not(t_59, y5);
not(t_60, t2);
or(e9, t_59, t_60);
and(f9, h0, x7);
not(t_61, v5);
not(t_62, u2);
or(g9, t_61, t_62);
and(h9, g0, w7);
not(t_63, c6);
not(t_64, v2);
or(i9, t_63, t_64);
and(j9, h6, f6, d6, b6);
and(k9, f0, v7);
not(t_65, a6);
not(t_66, w2);
or(l9, t_65, t_66);
and(m9, e0, u7);
not(t_67, g6);
not(t_68, x2);
or(n9, t_67, t_68);
and(o9, d0, t7);
not(t_69, e6);
not(t_70, y2);
or(p9, t_69, t_70);
and(q9, c0, s7);
and(r9, b0, r7);
not(t_71, v0);
not(t_72, a0);
not(t_73, p8);
or(s9, t_71, t_72, t_73);
and(t9, p8, a0, v0);
not(t_74, v0);
not(t_75, a0);
not(t_76, p8);
or(u9, t_74, t_75, t_76);
and(v9, p8, a0, v0);
not(t_77, a0);
not(t_78, p8);
or(w9, t_77, t_78);
and(x9, p8, a0);
and(y9, a3, e8);
and(z9, z, e8);
and(a10, n, o8);
not(b10, m6);
and(c10, d3, p6);
not(t_79, p6);
not(t_80, d3);
or(d10, t_79, t_80);
not(t_81, u6);
not(t_82, n6);
or(e10, t_81, t_82);
not(f10, n6);
not(t_83, t6);
not(t_84, o6);
or(g10, t_83, t_84);
not(h10, o6);
and(i10, q6, l8);
and(j10, g3, n8);
not(k10, r6);
not(l10, v6);
not(t_85, s6);
not(t_86, k);
or(m10, t_85, t_86);
and(n10, k, s6);
not(o10, w6);
and(p10, j, k8);
not(t_87, b7);
not(t_88, u3);
or(q10, t_87, t_88);
not(r10, x6);
not(t_89, g7);
not(t_90, z6);
or(s10, t_89, t_90);
not(t10, z6);
not(t_91, f7);
not(t_92, a7);
or(u10, t_91, t_92);
not(v10, a7);
and(w10, c7, h8);
and(x10, x3, j8);
not(y10, d7);
and(z10, b4, j7);
not(t_93, i7);
not(t_94, h7);
or(a11, t_93, t_94);
not(b11, h7);
not(c11, j7);
and(d11, l4, e7);
not(e11, l7);
not(f11, m7);
not(g11, n7);
not(h11, n7);
not(i11, n7);
not(j11, o7);
not(k11, p7);
not(l11, p7);
not(m11, p7);
not(n11, p7);
not(t_95, q7);
not(t_96, z7);
or(o11, t_95, t_96);
and(p11, a8, r4);
and(q11, a8, r4);
and(r11, a8, r4);
and(s11, a8, r4);
and(t11, a8, r4);
and(u11, a8, r4);
and(v11, a8, r4);
and(w11, a8, r4);
not(t_97, s4);
not(t_98, q8);
or(x11, t_97, t_98);
not(y11, a8);
not(z11, a8);
not(a12, a8);
not(b12, a8);
not(c12, a8);
not(d12, a8);
not(e12, a8);
not(f12, a8);
not(t_99, q7);
not(t_100, t4);
or(g12, t_99, t_100);
not(t_101, t4);
not(t_102, q8);
or(h12, t_101, t_102);
not(i12, b8);
not(j12, b8);
not(k12, b8);
not(l12, b8);
not(m12, b8);
not(n12, b8);
not(o12, b8);
and(p12, z4, f8);
and(q12, a5, f8);
not(r12, g8);
not(s12, g8);
not(t12, g8);
not(u12, g8);
not(v12, g8);
not(w12, g8);
not(x12, g8);
not(y12, g8);
and(z12, c5, g8);
and(a13, c5, g8);
and(b13, c5, g8);
and(c13, c5, g8);
and(d13, c5, g8);
and(e13, c5, g8);
and(f13, c5, g8);
and(g13, c5, g8);
not(t_103, z7);
not(t_104, d5);
not(t_105, f5);
or(h13, t_103, t_104, t_105);
not(t_106, e5);
not(t_107, t8);
not(t_108, n5);
or(i13, t_106, t_107, t_108);
not(j13, r8);
not(t_109, q7);
not(t_110, e5);
not(t_111, f5);
not(t_112, n5);
or(k13, t_109, t_110, t_111, t_112);
not(l13, s8);
not(t_113, z7);
not(t_114, f5);
or(m13, t_113, t_114);
not(n13, x8);
not(o13, x8);
not(p13, x8);
not(q13, x8);
not(r13, x8);
not(s13, x8);
not(t13, x8);
not(u13, x8);
and(v13, a, b, d8);
and(w13, a, b, c8);
or(x13, u8, a);
and(y13, l5, k7);
not(z13, y8);
not(t_115, l6);
not(t_116, t8);
not(t_117, n5);
or(a14, t_115, t_116, t_117);
not(t_118, x0);
not(t_119, z8);
or(b14, t_118, t_119);
and(c14, z8, x0);
and(d14, o0, f12);
and(e14, n0, e12);
and(f14, m0, d12);
and(g14, m0, y12);
not(t_120, c9);
not(t_121, a9);
or(h14, t_120, t_121);
not(t_122, b9);
not(t_123, j9);
or(i14, t_122, t_123);
and(j14, j0, w11);
and(k14, i0, v11);
not(t_124, g9);
not(t_125, e9);
or(l14, t_124, t_125);
and(m14, h0, u11);
and(n14, x5, j13);
and(o14, g0, t11);
not(t_126, l9);
not(t_127, i9);
or(p14, t_126, t_127);
and(q14, f0, s11);
and(r14, e0, r11);
not(t_128, p9);
not(t_129, n9);
or(s14, t_128, t_129);
and(t14, d0, q11);
and(u14, c0, p11);
buf(v14, u9);
not(t_130, p12);
not(t_131, i6);
or(w14, t_130, t_131);
not(t_132, q12);
not(t_133, i6);
or(x14, t_132, t_133);
not(t_134, y9);
not(t_135, i6);
or(y14, t_134, t_135);
not(t_136, z9);
not(t_137, i6);
or(z14, t_136, t_137);
not(t_138, p12);
not(t_139, j6);
or(a15, t_138, t_139);
not(t_140, q12);
not(t_141, j6);
or(b15, t_140, t_141);
not(t_142, y9);
not(t_143, j6);
or(c15, t_142, t_143);
not(t_144, z9);
not(t_145, j6);
or(d15, t_144, t_145);
and(e15, v, a13);
and(f15, u, z12);
not(t_146, n);
not(t_147, x13);
and(g15, t_146, t_147);
and(h15, n, c12);
and(i15, n, x12);
not(t_148, k10);
not(t_149, m6);
or(j15, t_148, t_149);
not(t_150, m);
not(t_151, x13);
and(k15, t_150, t_151);
and(l15, m, b12);
and(m15, m, w12);
not(t_152, b10);
not(t_153, r6);
or(n15, t_152, t_153);
not(t_154, l);
not(t_155, x13);
and(o15, t_154, t_155);
and(p15, l, a12);
not(t_156, h10);
not(t_157, j3);
or(q15, t_156, t_157);
not(t_158, f10);
not(t_159, k3);
or(r15, t_158, t_159);
and(s15, m3, v12);
and(t15, m3, g13);
not(t_160, o10);
not(t_161, v6);
or(u15, t_160, t_161);
not(t_162, k);
not(t_163, x13);
and(v15, t_162, t_163);
and(w15, k, z11);
and(x15, q3, u12);
and(y15, q3, f13);
not(t_164, l10);
not(t_165, w6);
or(z15, t_164, t_165);
not(t_166, j);
not(t_167, x13);
and(a16, t_166, t_167);
and(b16, j, y11);
and(c16, j, e13);
and(d16, j, t12);
not(t_168, y10);
not(t_169, x6);
or(e16, t_168, t_169);
not(t_170, i);
not(t_171, x13);
and(f16, t_170, t_171);
and(g16, y3, s12);
and(h16, y3, d13);
not(t_172, r10);
not(t_173, d7);
or(i16, t_172, t_173);
not(t_174, h);
not(t_175, x13);
and(j16, t_174, t_175);
not(t_176, v10);
not(t_177, c4);
or(k16, t_176, t_177);
not(t_178, t10);
not(t_179, d4);
or(l16, t_178, t_179);
and(m16, f4, r12);
and(n16, f4, c13);
and(o16, c10, y6, k4, h);
not(t_180, g);
not(t_181, x13);
and(p16, t_180, t_181);
and(q16, g, b13);
not(t_182, b11);
not(t_183, j4);
or(r16, t_182, t_183);
and(s16, d11, m7);
not(t16, o11);
and(u16, o11, g12);
and(v16, h12, x11);
not(w16, x11);
and(x16, h12, x11);
not(y16, x11);
not(z16, x11);
and(a17, h12, x11);
not(b17, x11);
and(c17, h12, x11);
not(d17, g12);
not(e17, h12);
not(f17, h12);
not(g17, h12);
not(h17, h12);
not(i17, h13);
not(j17, h13);
not(k17, h13);
not(l17, h13);
not(m17, i13);
not(n17, i13);
and(o17, i13, r8);
buf(p17, k13);
buf(q17, k13);
and(r17, s8, i13);
not(s17, m13);
not(t17, m13);
not(u17, m13);
not(v17, m13);
and(w17, x8, x13);
and(x17, x8, x13);
and(y17, x8, x13);
and(z17, x8, x13);
and(a18, x8, x13);
and(b18, x8, x13);
and(c18, x8, x13);
and(d18, x8, x13);
buf(e18, v13);
not(f18, v13);
buf(g18, w13);
not(h18, w13);
not(i18, y13);
not(j18, y13);
not(k18, y13);
not(l18, y13);
not(m18, y13);
not(n18, y13);
not(o18, y13);
not(p18, y13);
buf(q18, a14);
buf(r18, a14);
and(s18, h18, l0, n7);
and(t18, h18, l0, n7);
and(u18, h18, l0, n7);
and(v18, h18, l0, o7);
and(w18, f18, l0, p7);
and(x18, f18, l0, p7);
and(y18, f18, l0, p7);
and(z18, f18, l0, p7);
and(a19, h18, k0, i11);
not(b19, h14);
and(c19, i14, o17);
and(d19, h18, j0, h11);
and(e19, h18, i0, g11);
or(f19, j14, d9, d14);
not(g19, l14);
and(h19, h18, h0, j11);
or(i19, k14, f9, e14);
and(j19, f18, g0, n11);
or(k19, m14, h9, f14);
buf(l19, p14);
buf(m19, p14);
and(n19, f18, f0, m11);
or(o19, o14, k9, h15);
and(p19, f18, e0, l11);
or(q19, q14, m9, l15);
buf(r19, s14);
buf(s19, s14);
and(t19, f18, d0, k11);
or(u19, r14, o9, p15);
or(v19, t14, q9, w15);
or(w19, u14, r9, b16);
not(x19, v14);
buf(y19, w14);
buf(z19, w14);
buf(a20, x14);
buf(b20, x14);
buf(c20, y14);
buf(d20, y14);
buf(e20, z14);
buf(f20, z14);
buf(g20, a15);
buf(h20, a15);
buf(i20, b15);
buf(j20, b15);
buf(k20, c15);
buf(l20, c15);
buf(m20, d15);
buf(n20, d15);
and(o20, n, v8, d18);
or(p20, t15, g14, a10);
not(t_184, n15);
not(t_185, j15);
or(q20, t_184, t_185);
and(r20, d10, b17);
and(s20, d3, a17);
and(t20, m, v8, c18);
not(t_186, r15);
not(t_187, e10);
or(u20, t_186, t_187);
not(t_188, q15);
not(t_189, g10);
or(v20, t_188, t_189);
or(w20, h16, s15, i10);
or(x20, y15, i15, j10);
and(y20, h3, c17);
and(z20, l, v8, b18);
not(t_190, z15);
not(t_191, u15);
or(a21, t_190, t_191);
and(b21, n3, x16);
and(c21, k, v8, a18);
and(d21, m10, z16);
and(e21, r3, v16);
and(f21, j, w8, z17);
or(g21, n16, x15, p10);
not(t_192, i16);
not(t_193, e16);
or(h21, t_192, t_193);
and(i21, i, w8, y17);
not(t_194, l16);
not(t_195, s10);
or(j21, t_194, t_195);
not(t_196, k16);
not(t_197, u10);
or(k21, t_196, t_197);
or(l21, f15, m16, w10);
or(m21, q16, d16, x10);
and(n21, h, w8, x17);
not(t_198, r16);
not(t_199, a11);
or(o21, t_198, t_199);
and(p21, g, w8, w17);
and(q21, k4, u16);
and(r21, d11, m17);
and(s21, o16, l7);
and(t21, r18, h13);
and(u21, r18, h13);
and(v21, r18, h13);
and(w21, r18, h13);
not(x21, p17);
not(y21, p17);
not(z21, p17);
not(a22, p17);
not(b22, p17);
not(c22, p17);
not(d22, p17);
not(e22, p17);
not(f22, q17);
and(g22, q18, m13);
and(h22, q18, m13);
and(i22, q18, m13);
and(j22, q18, m13);
and(k22, y13, p17);
and(l22, y13, p17);
and(m22, y13, p17);
and(n22, y13, p17);
and(o22, y13, p17);
and(p22, y13, p17);
and(q22, y13, p17);
and(r22, y13, p17);
and(s22, q17, y8);
not(t22, q18);
not(u22, q18);
not(v22, q18);
not(w22, q18);
not(x22, r18);
not(y22, r18);
not(z22, r18);
not(a23, r18);
not(t_200, g19);
not(t_201, h14);
or(b23, t_200, t_201);
not(t_202, b19);
not(t_203, l14);
or(c23, t_202, t_203);
or(d23, c19, n14, r21);
not(t_204, r21);
not(t_205, n14);
not(t_206, c19);
and(e23, t_204, t_205, t_206);
not(f23, l19);
not(g23, m19);
not(h23, r19);
not(i23, s19);
not(j23, y19);
not(k23, y19);
not(l23, y19);
not(m23, y19);
not(n23, y19);
not(o23, y19);
not(p23, y19);
not(q23, y19);
not(r23, z19);
not(s23, z19);
not(t23, z19);
not(u23, z19);
not(v23, z19);
not(w23, z19);
not(x23, z19);
not(y23, z19);
not(z23, a20);
not(a24, a20);
not(b24, a20);
not(c24, a20);
not(d24, a20);
not(e24, a20);
not(f24, a20);
not(g24, a20);
not(h24, b20);
not(i24, b20);
not(j24, b20);
not(k24, b20);
not(l24, b20);
not(m24, b20);
not(n24, b20);
not(o24, b20);
not(p24, c20);
not(q24, c20);
not(r24, c20);
not(s24, c20);
not(t24, c20);
not(u24, c20);
not(v24, c20);
not(w24, c20);
not(x24, d20);
not(y24, d20);
not(z24, d20);
not(a25, d20);
not(b25, d20);
not(c25, d20);
not(d25, d20);
not(e25, d20);
not(f25, e20);
not(g25, e20);
not(h25, e20);
not(i25, e20);
not(j25, e20);
not(k25, e20);
not(l25, e20);
not(m25, e20);
not(n25, f20);
not(o25, f20);
not(p25, f20);
not(q25, f20);
not(r25, f20);
not(s25, f20);
not(t25, f20);
not(u25, f20);
not(v25, g20);
not(w25, g20);
not(x25, g20);
not(y25, g20);
not(z25, g20);
not(a26, g20);
not(b26, g20);
not(c26, g20);
not(d26, h20);
not(e26, h20);
not(f26, h20);
not(g26, h20);
not(h26, h20);
not(i26, h20);
not(j26, h20);
not(k26, h20);
not(l26, i20);
not(m26, i20);
not(n26, i20);
not(o26, i20);
not(p26, i20);
not(q26, i20);
not(r26, i20);
not(s26, i20);
not(t26, j20);
not(u26, j20);
not(v26, j20);
not(w26, j20);
not(x26, j20);
not(y26, j20);
not(z26, j20);
not(a27, j20);
not(b27, k20);
not(c27, k20);
not(d27, k20);
not(e27, k20);
not(f27, k20);
not(g27, k20);
not(h27, k20);
not(i27, k20);
not(j27, l20);
not(k27, l20);
not(l27, l20);
not(m27, l20);
not(n27, l20);
not(o27, l20);
not(p27, l20);
not(q27, l20);
not(r27, m20);
not(s27, m20);
not(t27, m20);
not(u27, m20);
not(v27, m20);
not(w27, m20);
not(x27, m20);
not(y27, m20);
not(z27, n20);
not(a28, n20);
not(b28, n20);
not(c28, n20);
not(d28, n20);
not(e28, n20);
not(f28, n20);
not(g28, n20);
not(h28, q20);
and(i28, c10, s22);
and(j28, e3, u20);
not(k28, v20);
not(l28, a21);
not(m28, h21);
and(n28, u3, j22);
and(o28, j21, v3, c11);
not(p28, k21);
and(q28, a4, i22);
not(r28, o21);
and(s28, g4, h22);
and(t28, k4, g22);
and(u28, d11, f22);
and(v28, l21, n13);
and(w28, m21, p13);
and(x28, g21, q13);
and(y28, w20, r13);
and(z28, x20, t13);
and(a29, p20, u13);
and(b29, e18, w19);
and(c29, e18, v19);
and(d29, e18, u19);
and(e29, e18, q19);
and(f29, g18, o19);
and(g29, g18, k19);
and(h29, g18, i19);
and(i29, g18, f19);
and(j29, t0, k26);
and(k29, s0, u25);
and(l29, s0, j26);
and(m29, r0, e25);
and(n29, r0, t25);
and(o29, r0, i26);
and(p29, q0, g28);
and(q29, q0, d25);
and(r29, q0, s25);
and(s29, q0, h26);
and(t29, p0, q27);
and(u29, p0, f28);
and(v29, p0, c25);
and(w29, p0, r25);
and(x29, p0, g26);
and(y29, o0, o24);
and(z29, o0, p27);
and(a30, o0, e28);
and(b30, o0, b25);
and(c30, o0, q25);
and(d30, o0, f26);
and(e30, n0, y23);
and(f30, n0, n24);
and(g30, n0, o27);
and(h30, n0, d28);
and(i30, n0, a25);
and(j30, n0, p25);
and(k30, n0, e26);
and(l30, m0, a27);
and(m30, m0, x23);
and(n30, m0, m24);
and(o30, m0, n27);
and(p30, m0, c28);
and(q30, m0, z24);
and(r30, m0, o25);
and(s30, m0, d26);
or(t30, i29, s18, a19);
or(u30, h29, t18, d19);
or(v30, g29, u18, e19);
or(w30, f29, v18, h19);
or(x30, e29, w18, j19);
or(y30, d29, x18, n19);
or(z30, c29, y18, p19);
or(a31, b29, z18, t19);
not(t_207, c23);
not(t_208, b23);
or(b31, t_207, t_208);
not(c31, e23);
not(t_209, h23);
not(t_210, l19);
or(d31, t_209, t_210);
not(t_211, i23);
not(t_212, m19);
or(e31, t_211, t_212);
not(t_213, f23);
not(t_214, r19);
or(f31, t_213, t_214);
not(t_215, g23);
not(t_216, s19);
or(g31, t_215, t_216);
and(h31, v, c26);
and(i31, v, l25);
and(j31, v, u24);
and(k31, v, v27);
and(l31, v, e27);
and(m31, v, b24);
and(n31, v, k23);
and(o31, v, l26);
and(p31, u, b26);
and(q31, u, k25);
and(r31, u, t24);
and(s31, u, u27);
and(t31, u, d27);
and(u31, u, a24);
and(v31, u, j23);
and(w31, t, a26);
and(x31, t, j25);
and(y31, t, s24);
and(z31, t, t27);
and(a32, t, c27);
and(b32, t, z23);
and(c32, s, z25);
and(d32, s, i25);
and(e32, s, r24);
and(f32, s, s27);
and(g32, s, b27);
and(h32, r, y25);
and(i32, r, h25);
and(j32, r, q24);
and(k32, r, r27);
and(l32, q, x25);
and(m32, q, g25);
and(n32, q, p24);
and(o32, p, w25);
and(p32, p, f25);
and(q32, o, v25);
or(r32, o20, g15, a29);
not(t_217, a29);
not(t_218, g15);
not(t_219, o20);
and(s32, t_217, t_218, t_219);
not(t_220, l28);
not(t_221, q20);
or(t32, t_220, t_221);
and(u32, e3, n25);
and(v32, e3, y24);
and(w32, e3, b28);
and(x32, e3, m27);
and(y32, e3, l24);
and(z32, e3, w23);
and(a33, e3, z26);
or(b33, t20, k15, z28);
not(t_222, z28);
not(t_223, k15);
not(t_224, t20);
and(c33, t_222, t_223, t_224);
and(d33, i3, s26);
and(e33, i3, x24);
and(f33, i3, a28);
and(g33, i3, l27);
and(h33, i3, k24);
and(i33, i3, v23);
and(j33, i3, y26);
not(t_225, h28);
not(t_226, a21);
or(k33, t_225, t_226);
and(l33, o3, r26);
and(m33, o3, q23);
and(n33, o3, z27);
and(o33, o3, k27);
and(p33, o3, j24);
and(q33, o3, u23);
and(r33, o3, x26);
or(s33, c21, v15, y28);
not(t_227, y28);
not(t_228, v15);
not(t_229, c21);
and(t33, t_227, t_228, t_229);
and(u33, s3, q26);
and(v33, s3, p23);
and(w33, s3, g24);
and(x33, s3, j27);
and(y33, s3, i24);
and(z33, s3, t23);
and(a34, s3, w26);
or(b34, f21, a16, x28);
not(t_230, x28);
not(t_231, a16);
not(t_232, f21);
and(c34, t_230, t_231, t_232);
and(d34, t3, p26);
and(e34, t3, o23);
and(f34, t3, f24);
and(g34, t3, i27);
and(h34, t3, h24);
and(i34, t3, s23);
and(j34, t3, v26);
not(t_233, r28);
not(t_234, h21);
or(k34, t_233, t_234);
or(l34, i21, f16, w28);
not(t_235, w28);
not(t_236, f16);
not(t_237, i21);
and(m34, t_235, t_236, t_237);
and(n34, z3, o26);
and(o34, z3, n23);
and(p34, z3, e24);
and(q34, z3, h27);
and(r34, z3, y27);
and(s34, z3, r23);
and(t34, z3, u26);
or(u34, z10, o28);
not(t_238, m28);
not(t_239, o21);
or(v34, t_238, t_239);
and(w34, h4, n26);
and(x34, h4, m23);
and(y34, h4, d24);
and(z34, h4, g27);
and(a35, h4, x27);
and(b35, h4, w24);
and(c35, h4, t26);
or(d35, p21, p16, v28);
not(t_240, v28);
not(t_241, p16);
not(t_242, p21);
and(e35, t_240, t_241, t_242);
and(f35, l4, m26);
and(g35, l4, l23);
and(h35, l4, c24);
and(i35, l4, f27);
and(j35, l4, w27);
and(k35, l4, v24);
and(l35, l4, m25);
and(m35, p28, i8);
and(n35, k28, m8);
and(o35, j28, n17);
not(t_243, j29);
not(t_244, l30);
not(t_245, e30);
not(t_246, y29);
not(t_247, t29);
not(t_248, p29);
not(t_249, m29);
not(t_250, k29);
and(p35, t_243, t_244, t_245, t_246, t_247, t_248, t_249, t_250);
not(t_251, l29);
not(t_252, a33);
not(t_253, m30);
not(t_254, f30);
not(t_255, z29);
not(t_256, u29);
not(t_257, q29);
not(t_258, n29);
and(q35, t_251, t_252, t_253, t_254, t_255, t_256, t_257, t_258);
not(t_259, o29);
not(t_260, j33);
not(t_261, z32);
not(t_262, n30);
not(t_263, g30);
not(t_264, a30);
not(t_265, v29);
not(t_266, r29);
and(r35, t_259, t_260, t_261, t_262, t_263, t_264, t_265, t_266);
not(t_267, s29);
not(t_268, r33);
not(t_269, i33);
not(t_270, y32);
not(t_271, o30);
not(t_272, h30);
not(t_273, b30);
not(t_274, w29);
and(s35, t_267, t_268, t_269, t_270, t_271, t_272, t_273, t_274);
not(t_275, x29);
not(t_276, a34);
not(t_277, q33);
not(t_278, h33);
not(t_279, x32);
not(t_280, p30);
not(t_281, i30);
not(t_282, c30);
and(t35, t_275, t_276, t_277, t_278, t_279, t_280, t_281, t_282);
not(t_283, d30);
not(t_284, j34);
not(t_285, z33);
not(t_286, p33);
not(t_287, g33);
not(t_288, w32);
not(t_289, q30);
not(t_290, j30);
and(u35, t_283, t_284, t_285, t_286, t_287, t_288, t_289, t_290);
not(t_291, k30);
not(t_292, t34);
not(t_293, i34);
not(t_294, y33);
not(t_295, o33);
not(t_296, f33);
not(t_297, v32);
not(t_298, r30);
and(v35, t_291, t_292, t_293, t_294, t_295, t_296, t_297, t_298);
not(t_299, s30);
not(t_300, c35);
not(t_301, s34);
not(t_302, h34);
not(t_303, x33);
not(t_304, n33);
not(t_305, e33);
not(t_306, u32);
and(w35, t_299, t_300, t_301, t_302, t_303, t_304, t_305, t_306);
buf(x35, t30);
not(y35, t30);
not(z35, t30);
buf(a36, u30);
not(b36, u30);
not(c36, u30);
buf(d36, v30);
not(e36, v30);
not(f36, v30);
buf(g36, w30);
not(h36, w30);
not(i36, w30);
buf(j36, x30);
not(k36, x30);
buf(l36, y30);
not(m36, y30);
buf(n36, z30);
not(o36, z30);
buf(p36, a31);
not(q36, a31);
buf(r36, b31);
not(t_307, f31);
not(t_308, d31);
or(s36, t_307, t_308);
not(t_309, g31);
not(t_310, e31);
or(t36, t_309, t_310);
and(u36, t9, b33);
and(v36, t9, r32);
and(w36, v9, l34);
and(x36, v9, b34);
and(y36, v9, s33);
and(z36, x9, d35);
and(a37, w30, v30, u30, t30, k6);
not(t_311, h31);
not(t_312, d33);
not(t_313, m33);
not(t_314, w33);
not(t_315, g34);
not(t_316, r34);
not(t_317, b35);
not(t_318, l35);
and(b37, t_311, t_312, t_313, t_314, t_315, t_316, t_317, t_318);
not(t_319, p31);
not(t_320, l33);
not(t_321, v33);
not(t_322, f34);
not(t_323, q34);
not(t_324, a35);
not(t_325, k35);
not(t_326, i31);
and(c37, t_319, t_320, t_321, t_322, t_323, t_324, t_325, t_326);
not(t_327, w31);
not(t_328, u33);
not(t_329, e34);
not(t_330, p34);
not(t_331, z34);
not(t_332, j35);
not(t_333, j31);
not(t_334, q31);
and(d37, t_327, t_328, t_329, t_330, t_331, t_332, t_333, t_334);
not(t_335, c32);
not(t_336, d34);
not(t_337, o34);
not(t_338, y34);
not(t_339, i35);
not(t_340, k31);
not(t_341, r31);
not(t_342, x31);
and(e37, t_335, t_336, t_337, t_338, t_339, t_340, t_341, t_342);
not(t_343, h32);
not(t_344, n34);
not(t_345, x34);
not(t_346, h35);
not(t_347, l31);
not(t_348, s31);
not(t_349, y31);
not(t_350, d32);
and(f37, t_343, t_344, t_345, t_346, t_347, t_348, t_349, t_350);
not(t_351, l32);
not(t_352, w34);
not(t_353, g35);
not(t_354, m31);
not(t_355, t31);
not(t_356, z31);
not(t_357, e32);
not(t_358, i32);
and(g37, t_351, t_352, t_353, t_354, t_355, t_356, t_357, t_358);
not(t_359, o32);
not(t_360, f35);
not(t_361, n31);
not(t_362, u31);
not(t_363, a32);
not(t_364, f32);
not(t_365, j32);
not(t_366, m32);
and(h37, t_359, t_360, t_361, t_362, t_363, t_364, t_365, t_366);
not(t_367, q32);
not(t_368, o31);
not(t_369, v31);
not(t_370, b32);
not(t_371, g32);
not(t_372, k32);
not(t_373, n32);
not(t_374, p32);
and(i37, t_367, t_368, t_369, t_370, t_371, t_372, t_373, t_374);
or(j37, e15, g16, m35);
not(k37, s32);
not(t_375, k33);
not(t_376, t32);
or(l37, t_375, t_376);
not(m37, c33);
or(n37, c16, m15, n35);
not(o37, t33);
not(p37, c34);
not(t_377, v34);
not(t_378, k34);
or(q37, t_377, t_378);
not(r37, m34);
not(s37, e35);
and(t37, b31, e17);
and(u37, u34, l13);
buf(v37, r36);
buf(w37, r36);
not(x37, s36);
buf(y37, t36);
buf(z37, t36);
buf(a38, u36);
buf(b38, u36);
buf(c38, v36);
buf(d38, v36);
buf(e38, w36);
buf(f38, w36);
buf(g38, x36);
buf(h38, x36);
buf(i38, y36);
buf(j38, y36);
buf(k38, z36);
buf(l38, z36);
and(m38, z, s32, x35);
and(n38, z, c33, a36);
and(o38, z, t33, g36);
and(p38, z, c34, j36);
and(q38, z, m34, l36);
and(r38, z, e35, p36);
and(s38, y, s32, y35);
and(t38, y, c33, b36);
and(u38, y, t33, h36);
and(v38, y, c34, k36);
and(w38, y, m34, m36);
and(x38, y, e35, q36);
and(y38, i36, f36, c36, z35, c3);
and(z38, x, r32, y35);
and(a39, x, b33, b36);
and(b39, x, s33, h36);
and(c39, x, b34, k36);
and(d39, x, l34, m36);
and(e39, x, d35, q36);
and(f39, w, r32, x35);
and(g39, w, b33, a36);
and(h39, w, s33, g36);
and(i39, w, b34, j36);
and(j39, w, l34, l36);
and(k39, w, d35, p36);
buf(l39, l37);
buf(m39, q37);
buf(n39, q37);
and(o39, q37, f11);
and(p39, i37, t16);
or(q39, e21, w16, t37);
and(r39, w35, d17);
and(s39, l37, f17);
and(t39, h37, i12);
and(u39, v35, b8);
and(v39, g37, j12);
and(w39, u35, b8);
and(x39, f37, k12);
and(y39, t35, b8);
and(z39, e37, l12);
and(a40, s35, b8);
and(b40, d37, m12);
and(c40, r35, b8);
and(d40, c37, n12);
and(e40, q35, b8);
and(f40, b37, o12);
and(g40, p35, b8);
and(h40, j37, o13);
and(i40, n37, s13);
not(j40, v37);
not(k40, w37);
not(l40, y37);
not(m40, z37);
not(n40, a38);
not(o40, b38);
not(p40, c38);
not(q40, d38);
not(r40, e38);
not(s40, f38);
not(t40, g38);
not(u40, h38);
not(v40, i38);
not(w40, j38);
not(x40, k38);
not(y40, l38);
or(z40, y38, a37);
or(a41, z38, f39);
not(t_379, f39);
not(t_380, z38);
and(b41, t_379, t_380);
or(c41, a39, g39);
not(t_381, g39);
not(t_382, a39);
and(d41, t_381, t_382);
or(e41, b39, h39);
not(t_383, h39);
not(t_384, b39);
and(f41, t_383, t_384);
or(g41, c39, i39);
not(t_385, i39);
not(t_386, c39);
and(h41, t_385, t_386);
or(i41, d39, j39);
not(t_387, j39);
not(t_388, d39);
and(j41, t_387, t_388);
or(k41, e39, k39);
not(t_389, k39);
not(t_390, e39);
and(l41, t_389, t_390);
or(m41, k37, m38, s38);
buf(n41, l39);
buf(o41, l39);
or(p41, m37, n38, t38);
or(q41, z20, o15, i40);
not(t_391, i40);
not(t_392, o15);
not(t_393, z20);
and(r41, t_391, t_392, t_393);
or(s41, o37, o38, u38);
or(t41, p37, p38, v38);
not(u41, m39);
not(v41, n39);
or(w41, r37, q38, w38);
or(x41, n21, j16, h40);
not(t_394, h40);
not(t_395, j16);
not(t_396, n21);
and(y41, t_394, t_395, t_396);
or(z41, s37, r38, x38);
or(a42, q21, r39, p39);
and(b42, x37, e11);
not(t_397, o39);
not(t_398, s16);
and(c42, t_397, t_398);
or(d42, b21, y16, s39);
or(e42, u39, t39);
or(f42, w39, v39);
or(g42, y39, x39);
or(h42, a40, z39);
or(i42, c40, b40);
or(j42, e40, d40);
or(k42, g40, f40);
and(l42, q39, t21);
not(t_399, l40);
not(t_400, v37);
or(m42, t_399, t_400);
not(t_401, m40);
not(t_402, w37);
or(n42, t_401, t_402);
not(t_403, j40);
not(t_404, y37);
or(o42, t_403, t_404);
not(t_405, k40);
not(t_406, z37);
or(p42, t_405, t_406);
and(q42, c41, s9);
and(r42, a41, s9);
and(s42, t9, q41);
and(t42, i41, u9);
and(u42, g41, u9);
and(v42, z40, x19);
and(w42, x9, x41);
and(x42, z, r41, d36);
and(y42, z, y41, n36);
and(z42, y, r41, e36);
and(a43, y, y41, o36);
and(b43, b41, m41);
and(c43, d41, p41);
and(d43, x, q41, e36);
not(e43, e41);
and(f43, f41, s41);
and(g43, h41, t41);
and(h43, j41, w41);
and(i43, x, x41, o36);
not(j43, k41);
and(k43, l41, z41);
and(l43, w, q41, d36);
and(m43, w, x41, n36);
not(t_407, u41);
not(t_408, n41);
or(n43, t_407, t_408);
not(o43, n41);
not(t_409, v41);
not(t_410, o41);
or(p43, t_409, t_410);
not(q43, o41);
not(r43, r41);
not(s43, y41);
not(t_411, b42);
not(t_412, s21);
and(t43, t_411, t_412);
and(u43, c42, g17);
and(v43, d42, u21);
and(w43, a42, t22);
and(x43, e42, u22);
and(y43, f42, v22);
and(z43, g42, w22);
and(a44, h42, x22);
and(b44, i42, y22);
and(c44, j42, z22);
and(d44, k42, a23);
not(t_413, o42);
not(t_414, m42);
or(e44, t_413, t_414);
not(t_415, p42);
not(t_416, n42);
or(f44, t_415, t_416);
buf(g44, r42);
buf(h44, r42);
buf(i44, s42);
buf(j44, s42);
not(k44, t42);
buf(l44, u42);
buf(m44, w42);
buf(n44, w42);
or(o44, r43, x42, z42);
or(p44, s43, y42, a43);
buf(q44, b43);
buf(r44, c43);
or(s44, d43, l43);
not(t_417, l43);
not(t_418, d43);
and(t44, t_417, t_418);
buf(u44, f43);
buf(v44, g43);
buf(w44, h43);
or(x44, i43, m43);
not(t_419, m43);
not(t_420, i43);
and(y44, t_419, t_420);
buf(z44, k43);
or(a45, s20, d21, u43);
not(t_421, o43);
not(t_422, m39);
or(b45, t_421, t_422);
not(t_423, q43);
not(t_424, n39);
or(c45, t_423, t_424);
and(d45, t43, h17);
not(e45, h44);
not(f45, i44);
not(g45, j44);
and(h45, s44, u9);
and(i45, x44, w9);
not(j45, m44);
not(k45, n44);
and(l45, t44, o44);
and(m45, y44, p44);
buf(n45, q44);
buf(o45, q44);
buf(p45, r44);
buf(q45, r44);
not(t_425, s44);
not(t_426, f43);
or(r45, t_425, t_426);
buf(s45, u44);
buf(t45, u44);
buf(u45, v44);
buf(v45, v44);
buf(w45, w44);
buf(x45, w44);
not(t_427, x44);
not(t_428, k43);
or(y45, t_427, t_428);
buf(z45, z44);
buf(a46, z44);
not(t_429, b45);
not(t_430, n43);
or(b46, t_429, t_430);
not(t_431, c45);
not(t_432, p43);
or(c46, t_431, t_432);
or(d46, y20, r20, d45);
and(e46, a45, w21);
not(t_433, n40);
not(t_434, p45);
or(f46, t_433, t_434);
not(t_435, o40);
not(t_436, q45);
or(g46, t_435, t_436);
not(t_437, p40);
not(t_438, n45);
or(h46, t_437, t_438);
not(t_439, q40);
not(t_440, o45);
or(i46, t_439, t_440);
not(j46, h45);
not(t_441, r40);
not(t_442, w45);
or(k46, t_441, t_442);
not(t_443, s40);
not(t_444, x45);
or(l46, t_443, t_444);
not(t_445, t40);
not(t_446, u45);
or(m46, t_445, t_446);
not(t_447, u40);
not(t_448, v45);
or(n46, t_447, t_448);
not(t_449, v40);
not(t_450, s45);
or(o46, t_449, t_450);
not(t_451, w40);
not(t_452, t45);
or(p46, t_451, t_452);
not(q46, i45);
not(t_453, x40);
not(t_454, z45);
or(r46, t_453, t_454);
not(t_455, y40);
not(t_456, a46);
or(s46, t_455, t_456);
buf(t46, l45);
buf(u46, m45);
not(t_457, f43);
not(t_458, c43);
not(t_459, l45);
not(t_460, a41);
or(v46, t_457, t_458, t_459, t_460);
and(w46, f43, l45, c43, b43);
not(x46, n45);
not(y46, o45);
not(t_461, c41);
not(t_462, l45);
not(t_463, f43);
or(z46, t_461, t_462, t_463);
not(a47, p45);
not(b47, q45);
not(c47, s45);
not(d47, t45);
not(t_464, k43);
not(t_465, h43);
not(t_466, m45);
not(t_467, g41);
or(e47, t_464, t_465, t_466, t_467);
and(f47, k43, m45, h43, g43);
not(g47, u45);
not(h47, v45);
not(t_468, i41);
not(t_469, m45);
not(t_470, k43);
or(i47, t_468, t_469, t_470);
not(j47, w45);
not(k47, x45);
not(l47, z45);
not(m47, a46);
not(n47, b46);
not(o47, c46);
and(p47, d46, v21);
not(t_471, a47);
not(t_472, a38);
or(q47, t_471, t_472);
not(t_473, b47);
not(t_474, b38);
or(r47, t_473, t_474);
not(t_475, x46);
not(t_476, c38);
or(s47, t_475, t_476);
not(t_477, y46);
not(t_478, d38);
or(t47, t_477, t_478);
and(u47, w46, v14);
not(t_479, j47);
not(t_480, e38);
or(v47, t_479, t_480);
not(t_481, k47);
not(t_482, f38);
or(w47, t_481, t_482);
not(t_483, g47);
not(t_484, g38);
or(x47, t_483, t_484);
not(t_485, h47);
not(t_486, h38);
or(y47, t_485, t_486);
not(t_487, c47);
not(t_488, i38);
or(z47, t_487, t_488);
not(t_489, d47);
not(t_490, j38);
or(a48, t_489, t_490);
not(t_491, l47);
not(t_492, k38);
or(b48, t_491, t_492);
not(t_493, m47);
not(t_494, l38);
or(c48, t_493, t_494);
buf(d48, t46);
buf(e48, t46);
buf(f48, u46);
buf(g48, u46);
not(t_495, v46);
not(t_496, z46);
not(t_497, r45);
not(t_498, e43);
or(h48, t_495, t_496, t_497, t_498);
buf(i48, f47);
not(t_499, e47);
not(t_500, i47);
not(t_501, y45);
not(t_502, j43);
or(j48, t_499, t_500, t_501, t_502);
and(k48, h48, s9);
not(t_503, f45);
not(t_504, d48);
or(l48, t_503, t_504);
not(t_505, g45);
not(t_506, e48);
or(m48, t_505, t_506);
not(t_507, f46);
not(t_508, q47);
or(n48, t_507, t_508);
not(t_509, g46);
not(t_510, r47);
or(o48, t_509, t_510);
not(t_511, h46);
not(t_512, s47);
or(p48, t_511, t_512);
not(t_513, i46);
not(t_514, t47);
or(q48, t_513, t_514);
or(r48, u47, v42);
not(t_515, k46);
not(t_516, v47);
or(s48, t_515, t_516);
not(t_517, l46);
not(t_518, w47);
or(t48, t_517, t_518);
not(t_519, m46);
not(t_520, x47);
or(u48, t_519, t_520);
not(t_521, n46);
not(t_522, y47);
or(v48, t_521, t_522);
not(t_523, o46);
not(t_524, z47);
or(w48, t_523, t_524);
not(t_525, p46);
not(t_526, a48);
or(x48, t_525, t_526);
not(t_527, r46);
not(t_528, b48);
or(y48, t_527, t_528);
not(t_529, s46);
not(t_530, c48);
or(z48, t_529, t_530);
not(t_531, j45);
not(t_532, f48);
or(a49, t_531, t_532);
not(t_533, k45);
not(t_534, g48);
or(b49, t_533, t_534);
not(c49, d48);
not(d49, e48);
not(e49, f48);
not(f49, g48);
not(t_535, h48);
not(t_536, f47);
or(g49, t_535, t_536);
not(h49, j48);
and(i49, u0, p48);
and(j49, u0, r48);
and(k49, n48, g44);
buf(l49, k48);
buf(m49, k48);
not(t_537, c49);
not(t_538, i44);
or(n49, t_537, t_538);
not(t_539, d49);
not(t_540, j44);
or(o49, t_539, t_540);
buf(p49, n48);
not(q49, o48);
buf(r49, p48);
not(s49, q48);
buf(t49, r48);
buf(u49, s48);
buf(v49, s48);
not(w49, t48);
buf(x49, u48);
buf(y49, u48);
not(z49, v48);
not(a50, w48);
not(b50, x48);
not(c50, y48);
not(d50, z48);
not(t_541, e49);
not(t_542, m44);
or(e50, t_541, t_542);
not(t_543, f49);
not(t_544, n44);
or(f50, t_543, t_544);
and(g50, g49, h49);
buf(h50, i49);
buf(i50, i49);
not(j50, j49);
or(k50, k49, q42);
not(t_545, e45);
not(t_546, p49);
or(l50, t_545, t_546);
and(m50, l49, x49);
not(t_547, l49);
not(t_548, y49);
not(t_549, v49);
or(n50, t_547, t_548, t_549);
not(o50, l49);
buf(p50, l49);
not(q50, m49);
not(t_550, l48);
not(t_551, n49);
or(r50, t_550, t_551);
not(t_552, m48);
not(t_553, o49);
or(s50, t_552, t_553);
and(t50, r49, n48);
not(u50, p49);
buf(v50, r49);
not(t_554, l44);
not(t_555, v49);
or(w50, t_554, t_555);
and(x50, t49, y49, v49);
and(y50, t49, x49);
buf(z50, v49);
buf(a51, x49);
not(t_556, a49);
not(t_557, e50);
or(b51, t_556, t_557);
not(t_558, b49);
not(t_559, f50);
or(c51, t_558, t_559);
and(d51, l49, i48);
and(e51, t49, i48);
and(f51, b50, i17);
and(g51, q49, k17);
and(h51, s49, l17);
and(i51, d50, s17);
and(j51, w49, u17);
and(k51, z49, v17);
and(l51, u0, r48, o50);
not(t_560, q5);
not(t_561, v50);
or(m51, t_560, t_561);
not(n51, h50);
not(o51, i50);
and(p51, u0, t50);
and(q51, u0, y50);
and(r51, u0, x50);
not(t_562, q42);
not(t_563, r50);
or(s51, t_562, t_563);
buf(t51, k50);
buf(u51, k50);
not(t_564, g44);
not(t_565, n48);
not(t_566, r50);
or(v51, t_564, t_565, t_566);
not(t_567, u50);
not(t_568, h44);
or(w51, t_567, t_568);
not(t_569, q50);
not(t_570, a51);
or(x51, t_569, t_570);
buf(y51, r50);
not(z51, s50);
and(a52, r49, n48, r50);
not(b52, v50);
not(t_571, n50);
not(t_572, w50);
not(t_573, k44);
or(c52, t_571, t_572, t_573);
or(d52, m50, u42);
not(e52, z50);
not(f52, a51);
buf(g52, b51);
buf(h52, b51);
not(i52, c51);
buf(j52, e51);
or(k52, d51, j48);
not(t_574, z43);
not(t_575, k51);
not(t_576, n28);
and(l52, t_574, t_575, t_576);
not(t_577, y43);
not(t_578, j51);
not(t_579, q28);
and(m52, t_577, t_578, t_579);
not(t_580, w43);
not(t_581, i51);
not(t_582, t28);
and(n52, t_580, t_581, t_582);
not(t_583, a44);
not(t_584, f51);
not(t_585, l42);
and(o52, t_583, t_584, t_585);
not(t_586, c44);
not(t_587, g51);
not(t_588, p47);
and(p52, t_586, t_587, t_588);
not(t_589, d44);
not(t_590, h51);
not(t_591, e46);
and(q52, t_589, t_590, t_591);
not(t_592, b52);
not(t_593, p2);
or(r52, t_592, t_593);
not(s52, p51);
and(t52, u0, a52);
buf(u52, q51);
buf(v52, q51);
not(w52, r51);
and(x52, k50, u51);
not(y52, t51);
not(z52, u51);
not(t_594, w51);
not(t_595, l50);
or(a53, t_594, t_595);
not(t_596, l49);
not(t_597, y49);
not(t_598, u49);
not(t_599, h52);
or(b53, t_596, t_597, t_598, t_599);
or(c53, p50, l51);
not(t_600, l51);
not(t_601, p50);
and(d53, t_600, t_601);
not(t_602, f52);
not(t_603, m49);
or(e53, t_602, t_603);
not(f53, y51);
not(t_604, t42);
not(t_605, h52);
or(g53, t_604, t_605);
not(h53, c52);
not(t_606, l44);
not(t_607, u49);
not(t_608, h52);
or(i53, t_606, t_607, t_608);
not(t_609, e52);
not(t_610, d52);
or(j53, t_609, t_610);
not(k53, d52);
not(t_611, v51);
not(t_612, s51);
not(t_613, j46);
or(l53, t_611, t_612, t_613);
and(m53, t49, h52, v49, y49);
not(n53, g52);
not(o53, j52);
buf(p53, k52);
buf(q53, k52);
and(r53, z51, j17);
and(s53, i52, t17);
and(t53, n52, k22);
and(u53, m52, m22);
and(v53, l52, n22);
and(w53, o52, o22);
and(x53, p52, q22);
and(y53, q52, r22);
and(z53, u0, t50, z52);
not(t_614, r52);
not(t_615, m51);
or(a54, t_614, t_615);
buf(b54, t52);
buf(c54, t52);
not(d54, u52);
not(e54, v52);
and(f54, u0, m53);
not(t_616, f53);
not(t_617, t51);
or(g54, t_616, t_617);
buf(h54, a53);
buf(i54, a53);
buf(j54, d53);
not(t_618, e53);
not(t_619, x51);
or(k54, t_618, t_619);
not(t_620, y52);
not(t_621, y51);
or(l54, t_620, t_621);
not(t_622, n53);
not(t_623, c52);
or(m54, t_622, t_623);
not(n54, l53);
buf(o54, m53);
not(t_624, k53);
not(t_625, z50);
or(p54, t_624, t_625);
not(t_626, a50);
not(t_627, l53);
or(q54, t_626, t_627);
not(t_628, b53);
not(t_629, i53);
not(t_630, g53);
not(t_631, q46);
or(r54, t_628, t_629, t_630, t_631);
not(t_632, h53);
not(t_633, g52);
or(s54, t_632, t_633);
not(t54, p53);
not(u54, q53);
and(v54, k52, q53);
not(t_634, x43);
not(t_635, s53);
not(t_636, s28);
and(w54, t_634, t_635, t_636);
not(t_637, b44);
not(t_638, r53);
not(t_639, v43);
and(x54, t_637, t_638, t_639);
and(y54, c53, z13);
and(z54, u0, e51, u54);
not(t_640, n51);
not(t_641, h54);
or(a55, t_640, t_641);
not(t_642, o51);
not(t_643, i54);
or(b55, t_642, t_643);
not(c55, b54);
not(d55, c54);
not(t_644, j50);
not(t_645, k54);
or(e55, t_644, t_645);
buf(f55, f54);
buf(g55, f54);
not(t_646, g54);
not(t_647, l54);
or(h55, t_646, t_647);
not(i55, h54);
not(j55, i54);
buf(k55, j54);
not(l55, k54);
not(t_648, m54);
not(t_649, s54);
or(m55, t_648, t_649);
not(t_650, j53);
not(t_651, p54);
or(n55, t_650, t_651);
not(o55, o54);
not(t_652, n54);
not(t_653, w48);
or(p55, t_652, t_653);
buf(q55, r54);
buf(r55, r54);
not(t_654, o53);
not(t_655, o54);
or(s55, t_654, t_655);
or(t55, i28, y54, u28);
not(t_656, u28);
not(t_657, y54);
not(t_658, i28);
and(u55, t_656, t_657, t_658);
and(v55, a54, e22);
and(w55, w54, l22);
and(x55, x54, p22);
and(y55, a54, p18);
not(t_659, i55);
not(t_660, h50);
or(z55, t_659, t_660);
not(t_661, j55);
not(t_662, i50);
or(a56, t_661, t_662);
not(t_663, s52);
not(t_664, h55);
or(b56, t_663, t_664);
not(t_665, l55);
not(t_666, j49);
or(c56, t_665, t_666);
not(t_667, w52);
not(t_668, m55);
or(d56, t_667, t_668);
not(e56, f55);
not(f56, g55);
not(g56, h55);
not(h56, k55);
not(i56, m55);
buf(j56, n55);
buf(k56, n55);
not(t_669, q54);
not(t_670, p55);
or(l56, t_669, t_670);
not(m56, q55);
not(n56, r55);
not(t_671, c50);
not(t_672, r55);
or(o56, t_671, t_672);
not(t_673, o55);
not(t_674, j52);
or(p56, t_673, t_674);
not(t_675, t54);
not(t_676, q55);
or(q56, t_675, t_676);
not(t_677, z54);
not(t_678, v54);
and(r56, t_677, t_678);
not(s56, u55);
or(t56, y53, v55, y55);
not(t_679, y55);
not(t_680, v55);
not(t_681, y53);
and(u56, t_679, t_680, t_681);
not(t_682, a55);
not(t_683, z55);
or(v56, t_682, t_683);
not(t_684, b55);
not(t_685, a56);
or(w56, t_684, t_685);
not(t_686, g56);
not(t_687, p51);
or(x56, t_686, t_687);
not(t_688, e55);
not(t_689, c56);
or(y56, t_688, t_689);
not(t_690, d54);
not(t_691, j56);
or(z56, t_690, t_691);
not(t_692, e54);
not(t_693, k56);
or(a57, t_692, t_693);
not(t_694, i56);
not(t_695, r51);
or(b57, t_694, t_695);
not(c57, j56);
not(d57, k56);
buf(e57, l56);
buf(f57, l56);
not(t_696, n56);
not(t_697, y48);
or(g57, t_696, t_697);
not(t_698, p56);
not(t_699, s55);
or(h57, t_698, t_699);
not(t_700, m56);
not(t_701, p53);
or(i57, t_700, t_701);
buf(j57, r56);
buf(k57, t56);
not(l57, u56);
not(m57, w56);
not(t_702, b56);
not(t_703, x56);
or(n57, t_702, t_703);
not(t_704, c55);
not(t_705, e57);
or(o57, t_704, t_705);
not(t_706, d55);
not(t_707, f57);
or(p57, t_706, t_707);
not(t_708, c57);
not(t_709, u52);
or(q57, t_708, t_709);
not(t_710, d57);
not(t_711, v52);
or(r57, t_710, t_711);
not(t_712, d56);
not(t_713, b57);
or(s57, t_712, t_713);
and(t57, u0, h57);
and(u57, v56, d53);
not(v57, e57);
not(w57, f57);
not(t_714, o56);
not(t_715, g57);
or(x57, t_714, t_715);
not(t_716, q56);
not(t_717, i57);
or(y57, t_716, t_717);
buf(z57, j57);
and(a58, y56, a22);
and(b58, y56, l18);
and(c58, v56, o18);
not(d58, k57);
not(e58, m57);
buf(f58, n57);
not(t_718, v57);
not(t_719, b54);
or(g58, t_718, t_719);
not(t_720, w57);
not(t_721, c54);
or(h58, t_720, t_721);
not(t_722, z56);
not(t_723, q57);
or(i58, t_722, t_723);
not(t_724, a57);
not(t_725, r57);
or(j58, t_724, t_725);
buf(k58, s57);
not(l58, t57);
not(t_726, h56);
not(t_727, m57);
or(m58, t_726, t_727);
not(n58, u57);
buf(o58, x57);
buf(p58, x57);
not(q58, y57);
not(r58, z57);
and(s58, s57, j18);
or(t58, v53, a58, b58);
not(t_728, b58);
not(t_729, a58);
not(t_730, v53);
and(u58, t_728, t_729, t_730);
and(v58, n57, n18);
not(t_731, n58);
not(t_732, f58);
or(w58, t_731, t_732);
not(x58, f58);
not(t_733, o57);
not(t_734, g58);
or(y58, t_733, t_734);
not(t_735, p57);
not(t_736, h58);
or(z58, t_735, t_736);
not(a59, j58);
not(b59, k58);
not(t_737, e56);
not(t_738, o58);
or(c59, t_737, t_738);
not(t_739, f56);
not(t_740, p58);
or(d59, t_739, t_740);
not(t_741, q58);
not(t_742, t57);
or(e59, t_741, t_742);
not(t_743, e58);
not(t_744, k55);
or(f59, t_743, t_744);
not(g59, o58);
not(h59, p58);
not(t_745, l58);
not(t_746, y57);
or(i59, t_745, t_746);
and(j59, i58, r56);
and(k59, i58, k18);
buf(l59, t58);
buf(m59, t58);
not(n59, u58);
not(o59, z58);
not(p59, a59);
not(t_747, b59);
not(t_748, j59);
or(q59, t_747, t_748);
not(t_749, g59);
not(t_750, f55);
or(r59, t_749, t_750);
not(t_751, h59);
not(t_752, g55);
or(s59, t_751, t_752);
not(t_753, i59);
not(t_754, e59);
or(t59, t_753, t_754);
and(u59, v56, n57, y58, j54);
not(t_755, m58);
not(t_756, f59);
or(v59, t_755, t_756);
not(t_757, x58);
not(t_758, u57);
or(w59, t_757, t_758);
not(t_759, r58);
not(t_760, a59);
or(x59, t_759, t_760);
not(y59, j59);
not(z59, l59);
not(a60, m59);
and(b60, y58, m18);
not(t_761, w58);
not(t_762, w59);
or(c60, t_761, t_762);
not(t_763, y59);
not(t_764, k58);
or(d60, t_763, t_764);
not(t_765, c59);
not(t_766, r59);
or(e60, t_765, t_766);
not(t_767, d59);
not(t_768, s59);
or(f60, t_767, t_768);
not(t_769, o59);
not(t_770, j54);
and(g60, t_769, t_770);
not(h60, v59);
not(t_771, p59);
not(t_772, z57);
or(i60, t_771, t_772);
and(j60, t59, r17);
not(t_773, d60);
not(t_774, q59);
or(k60, t_773, t_774);
not(l60, f60);
or(m60, u59, g60);
and(n60, i58, s57, e60, j57);
not(t_775, x59);
not(t_776, i60);
or(o60, t_775, t_776);
or(p60, j60, o35, u37);
not(t_777, u37);
not(t_778, o35);
not(t_779, j60);
and(q60, t_777, t_778, t_779);
and(r60, c60, c22);
and(s60, h60, d22);
and(t60, e60, i18);
not(t_780, l60);
not(t_781, j57);
and(u60, t_780, t_781);
not(v60, o60);
not(w60, q60);
and(x60, k60, y21);
and(y60, m60, b22);
or(z60, x55, r60, v58);
not(t_782, v58);
not(t_783, r60);
not(t_784, x55);
and(a61, t_782, t_783, t_784);
or(b61, x53, s60, c58);
not(t_785, c58);
not(t_786, s60);
not(t_787, x53);
and(c61, t_785, t_786, t_787);
or(d61, n60, u60);
and(e61, v60, z21);
or(n1, w55, x60, s58);
not(t_788, s58);
not(t_789, x60);
not(t_790, w55);
and(g61, t_788, t_789, t_790);
or(h61, w53, y60, b60);
not(t_791, b60);
not(t_792, y60);
not(t_793, w53);
and(i61, t_791, t_792, t_793);
buf(j61, z60);
not(k61, a61);
buf(l61, b61);
not(m61, c61);
and(n61, n1, o5);
and(o61, d61, x21);
buf(p61, n1);
or(q61, u53, e61, k59);
not(t_794, k59);
not(t_795, e61);
not(t_796, u53);
and(r61, t_794, t_795, t_796);
buf(s61, h61);
not(t61, i61);
not(u61, j61);
not(v61, l61);
not(t_797, d58);
not(t_798, l61);
or(w61, t_797, t_798);
and(x61, u56, c61, a61, i61);
buf(y61, n61);
buf(z61, n61);
or(o1, t53, o61, t60);
not(t_799, t60);
not(t_800, o61);
not(t_801, t53);
and(b62, t_799, t_800, t_801);
not(c62, p61);
buf(d62, q61);
not(e62, r61);
not(t_802, u61);
not(t_803, s61);
or(f62, t_802, t_803);
not(g62, s61);
not(t_804, v61);
not(t_805, k57);
or(h62, t_804, t_805);
and(i62, o5, o1);
not(j62, y61);
not(k62, z61);
and(l62, g61, b62, p5);
buf(m62, o1);
buf(n62, d62);
buf(o62, d62);
and(p62, u58, r61, g61, b62);
not(t_806, g62);
not(t_807, j61);
or(q62, t_806, t_807);
not(t_808, h62);
not(t_809, w61);
or(r62, t_808, t_809);
buf(s62, i62);
buf(t62, i62);
not(u62, m62);
not(t_810, c62);
not(t_811, m62);
or(v62, t_810, t_811);
not(w62, n62);
not(x62, o62);
not(t_812, z59);
not(t_813, n62);
or(y62, t_812, t_813);
not(t_814, a60);
not(t_815, o62);
or(z62, t_814, t_815);
not(t_816, q62);
not(t_817, f62);
or(a63, t_816, t_817);
buf(b63, r62);
buf(c63, r62);
and(d63, x61, p62);
and(e63, x61, p62);
not(f63, s62);
not(g63, t62);
not(t_818, j62);
not(t_819, s62);
or(h63, t_818, t_819);
not(t_820, k62);
not(t_821, t62);
or(i63, t_820, t_821);
not(t_822, l62);
not(t_823, e63);
and(j63, t_822, t_823);
not(t_824, u62);
not(t_825, p61);
or(k63, t_824, t_825);
not(t_826, w62);
not(t_827, l59);
or(l63, t_826, t_827);
not(t_828, x62);
not(t_829, m59);
or(m63, t_828, t_829);
buf(n63, a63);
buf(o63, a63);
not(p63, b63);
not(q63, c63);
not(t_830, f63);
not(t_831, y61);
or(r63, t_830, t_831);
not(t_832, g63);
not(t_833, z61);
or(s63, t_832, t_833);
and(t63, a0, j63);
not(t_834, k63);
not(t_835, v62);
or(u63, t_834, t_835);
not(t_836, l63);
not(t_837, y62);
or(v63, t_836, t_837);
not(t_838, m63);
not(t_839, z62);
or(w63, t_838, t_839);
not(t_840, p63);
not(t_841, n63);
or(x63, t_840, t_841);
not(y63, n63);
not(t_842, q63);
not(t_843, o63);
or(z63, t_842, t_843);
not(a64, o63);
not(t_844, h63);
not(t_845, r63);
or(b64, t_844, t_845);
not(t_846, i63);
not(t_847, s63);
or(c64, t_846, t_847);
not(d64, u63);
buf(e64, v63);
not(f64, w63);
not(t_848, y63);
not(t_849, b63);
or(g64, t_848, t_849);
not(t_850, a64);
not(t_851, c63);
or(h64, t_850, t_851);
and(i64, f64, b64, b14);
and(j64, v63, b64, c14);
not(k64, c64);
not(t_852, d64);
not(t_853, e64);
or(l64, t_852, t_853);
not(m64, e64);
not(t_854, g64);
not(t_855, x63);
or(n64, t_854, t_855);
not(t_856, h64);
not(t_857, z63);
or(o64, t_856, t_857);
and(p64, v63, k64, b14);
and(q64, f64, k64, c14);
not(t_858, m64);
not(t_859, u63);
or(r64, t_858, t_859);
buf(s64, n64);
buf(t64, n64);
not(u64, o64);
or(v64, q64, i64, p64, j64);
not(t_860, l64);
not(t_861, r64);
or(w64, t_860, t_861);
not(x64, s64);
not(y64, t64);
buf(z64, u64);
buf(a65, u64);
buf(b65, v64);
buf(c65, v64);
buf(d65, w64);
buf(e65, w64);
not(f65, z64);
not(g65, a65);
not(t_862, f65);
not(t_863, b65);
or(h65, t_862, t_863);
not(i65, b65);
not(t_864, g65);
not(t_865, c65);
or(j65, t_864, t_865);
not(k65, c65);
not(l65, d65);
not(m65, e65);
not(t_866, x64);
not(t_867, d65);
or(n65, t_866, t_867);
not(t_868, y64);
not(t_869, e65);
or(o65, t_868, t_869);
not(t_870, l65);
not(t_871, s64);
or(p65, t_870, t_871);
not(t_872, m65);
not(t_873, t64);
or(q65, t_872, t_873);
not(t_874, i65);
not(t_875, z64);
or(r65, t_874, t_875);
not(t_876, k65);
not(t_877, a65);
or(s65, t_876, t_877);
not(t_878, h65);
not(t_879, r65);
or(t65, t_878, t_879);
not(t_880, j65);
not(t_881, s65);
or(u65, t_880, t_881);
not(t_882, p65);
not(t_883, n65);
or(v65, t_882, t_883);
not(t_884, q65);
not(t_885, o65);
or(w65, t_884, t_885);
endmodule
module top;
	parameter in_width = 50,
		patterns = 5000,
		step = 1;
	reg [1:in_width] in_mem[1:patterns];
	integer index;

	wire i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,
		i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,
		i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,
		i30,i31,i32,i33,i34,i35,i36,i37,i38,i39,
		i40,i41,i42,i43,i44,i45,i46,i47,i48,i49;

	assign {i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,
		i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,
		i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,
		i30,i31,i32,i33,i34,i35,i36,i37,i38,i39,
		i40,i41,i42,i43,i44,i45,i46,i47,i48,i49} = 
		$getpattern(in_mem[index]);

	initial $monitor($time,,o0,o1,o2,o3,o4,o5,o6,o7,o8,o9,
		o10,o11,o12,o13,o14,o15,o16,o17,o18,o19,
		o20,o21);
	initial
		begin
			$readmemb("patt.mem", in_mem);
			for(index = 1; index <= patterns; index = index + 1)
				#step;
		end

	foobar cct(o0,o1,o2,o3,o4,o5,o6,o7,o8,o9,
		o10,o11,o12,o13,o14,o15,o16,o17,o18,o19,
		o20,o21,i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,
		i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,
		i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,
		i30,i31,i32,i33,i34,i35,i36,i37,i38,i39,
		i40,i41,i42,i43,i44,i45,i46,i47,i48,i49);
endmodule