// IWLS benchmark module "ttt2" printed on Wed May 29 16:25:17 2002
module ttt2(a, b, c, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, \x , y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0);
input
  a,
  b,
  c,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  t,
  u,
  v,
  w,
  \x ,
  y;
output
  g0,
  h0,
  i0,
  j0,
  k0,
  l0,
  m0,
  z,
  n0,
  o0,
  p0,
  q0,
  r0,
  s0,
  t0,
  a0,
  b0,
  c0,
  d0,
  e0,
  f0;
wire
  \[26] ,
  \[27] ,
  \[28] ,
  j2,
  \[29] ,
  k2,
  \[10] ,
  \[45] ,
  \[11] ,
  \[12] ,
  \[13] ,
  \[48] ,
  o2,
  \[14] ,
  \[49] ,
  \[0] ,
  \[15] ,
  \[30] ,
  \[1] ,
  \[16] ,
  \[31] ,
  \[2] ,
  \[17] ,
  \[32] ,
  \[3] ,
  \[18] ,
  \[33] ,
  \[4] ,
  \[19] ,
  \[5] ,
  \[6] ,
  w1,
  w3,
  \[36] ,
  \[7] ,
  \[37] ,
  \[8] ,
  \[38] ,
  \[9] ,
  z1,
  \[39] ,
  a3,
  \[20] ,
  \[21] ,
  \[23] ,
  \[24] ,
  f3,
  \[25] ;
assign
  g0 = \[7] ,
  \[26]  = \[23]  | t,
  h0 = \[8] ,
  \[27]  = \[24]  | \[21] ,
  i0 = \[9] ,
  \[28]  = \[26]  | y,
  j0 = \[10] ,
  j2 = (v & u) | (~u & t),
  \[29]  = (~j2 & s) | (~y & ~v),
  k0 = \[11] ,
  k2 = (y & (~v & (~t & (~s & q)))) | \[49] ,
  \[10]  = (~w3 & (~o & ~a)) | (w3 & (o & ~a)),
  \[45]  = \[27]  | ~o,
  l0 = \[12] ,
  \[11]  = (~\[24]  & (\[21]  & ~f3)) | ((w3 & (~f3 & p)) | (~f3 & ~o)),
  m0 = \[13] ,
  \[12]  = (~\[30]  & (~\[10]  & (~q & ~a))) | ((\[30]  & (q & ~a)) | (\[10]  & q)),
  z = \[0] ,
  n0 = \[14] ,
  \[13]  = (~\[30]  & (~r & (q & (o & ~a)))) | ((~f3 & (r & (q & ~p))) | ((\[38]  & (~f3 & r)) | ((\[31]  & (\[6]  & r)) | ((~\[21]  & (p & ~a)) | (r & (~o & ~a)))))),
  \[48]  = ~j2 & t,
  o0 = \[15] ,
  o2 = (~z1 & (v & ~s)) | ((\[39]  & ~j) | (~\[23]  & t)),
  \[14]  = (~\[45]  & \[33] ) | (\[45]  & \[32] ),
  \[49]  = ~v & ~u,
  p0 = \[16] ,
  \[0]  = (j2 & (~w & e)) | ((\[49]  & ~w) | (~\[25]  & ~w)),
  \[15]  = (\[32]  & (~\[27]  & (j2 & (~\[10]  & ~t)))) | ((~\[27]  & (~\[26]  & (~\[10]  & ~a))) | ((\[27]  & (t & ~a)) | ((\[33]  & t) | (\[10]  & t)))),
  q0 = \[17] ,
  \[30]  = w3 | ~p,
  \[1]  = (\[37]  & (w & ~q)) | ((~w1 & (~w & v)) | (~w1 & ~q)),
  \[16]  = (\[32]  & (z1 & (~\[14]  & ~u))) | ((z1 & (~t & ~a)) | ((\[33]  & u) | (\[14]  & u))),
  r0 = \[18] ,
  \[31]  = ~\x  | ~o,
  \[2]  = (\[39]  & (~w & g)) | ((\[29]  & (~w & u)) | ((\[48]  & ~w) | ~\[37] )),
  \[17]  = (\[48]  & (\[32]  & ~\[14] )) | ((\[33]  & v) | ((\[16]  & v) | (\[14]  & v))),
  s0 = \[19] ,
  \[32]  = s & ~a,
  \[3]  = (\[25]  & (~k2 & (~j2 & ~w))) | ((\[25]  & (~k2 & (~w & h))) | ((w & ~q) | ~\[36] )),
  \[18]  = (\[33]  & (z1 & (y & (~v & ~t)))) | (\[36]  & (w & ~a)),
  t0 = \[20] ,
  \[33]  = ~s & ~a,
  \[4]  = (\[39]  & (~w & i)) | (~\[23]  & (j2 & ~w)),
  \[19]  = (~\x  & (b & ~a)) | (\x  & (~b & ~a)),
  \[5]  = (~o2 & (~w & v)) | (~o2 & (~w & ~u)),
  \[6]  = ~a & ~k,
  w1 = (j2 & ~f) | (\[49]  | (\[48]  | \[29] )),
  w3 = a3 & ~\x ,
  \[36]  = \[28]  | ~z1,
  \[7]  = (a3 & (~\[6]  & (~l & ~a))) | (\[6]  & l),
  \[37]  = \[28]  | ~u,
  \[8]  = (~m & (l & (k & ~a))) | ((m & (~l & ~a)) | (\[6]  & m)),
  \[38]  = ~n | (m | l),
  \[9]  = (~\[8]  & (~n & (m & ~a))) | ((\[8]  & n) | (\[6]  & n)),
  z1 = t | u,
  \[39]  = z1 & v,
  a0 = \[1] ,
  a3 = \[38]  | ~k,
  \[20]  = (~y & (c & ~a)) | (y & (~c & ~a)),
  b0 = \[2] ,
  \[21]  = ~r | q,
  c0 = \[3] ,
  d0 = \[4] ,
  \[23]  = v | ~s,
  e0 = \[5] ,
  \[24]  = w3 | p,
  f0 = \[6] ,
  f3 = (~\[31]  & ~\[21] ) | ((~\[31]  & p) | ((~p & ~o) | a)),
  \[25]  = z1 | ~s;
endmodule

