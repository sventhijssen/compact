// IWLS benchmark module "lal" printed on Wed May 29 16:09:11 2002
module lal(a, b, c, d, e, f, g, h, j, k, l, m, n, o, p, q, r, s, t, u, v, w, \x , y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0);
input
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  t,
  u,
  v,
  w,
  \x ,
  y,
  z,
  a0;
output
  k0,
  l0,
  m0,
  n0,
  o0,
  p0,
  q0,
  r0,
  s0,
  t0,
  b0,
  c0,
  d0,
  e0,
  f0,
  g0,
  h0,
  i0,
  j0;
wire
  \[13] ,
  \[14] ,
  \[15] ,
  \[16] ,
  \[17] ,
  p2,
  \[18] ,
  q1,
  \[19] ,
  \[0] ,
  \[1] ,
  t2,
  t3,
  \[3] ,
  d2,
  \[4] ,
  \[5] ,
  \[20] ,
  \[6] ,
  \[7] ,
  \[22] ,
  \[8] ,
  \[10] ,
  \[23] ,
  \[9] ,
  \[11] ,
  \[24] ,
  \[12] ;
assign
  k0 = \[9] ,
  \[13]  = (d2 & v) | (~\[22]  | q1),
  l0 = \[10] ,
  \[14]  = (\[22]  & w) | (~\[19]  | q1),
  m0 = \[11] ,
  \[15]  = (\[19]  & \x ) | (~\[24]  | q1),
  n0 = \[12] ,
  \[16]  = (\[24]  & y) | (t2 | q1),
  o0 = \[13] ,
  \[17]  = (~t2 & z) | ((t2 & ~z) | q1),
  p0 = \[14] ,
  p2 = w | v,
  \[18]  = (t2 & (\[17]  & ~a0)) | ((~t2 & a0) | ((~\[17]  & a0) | q1)),
  q0 = \[15] ,
  q1 = \[9]  | (q | h),
  \[19]  = p2 | d2,
  r0 = \[16] ,
  s0 = \[17] ,
  \[0]  = j & ~r,
  t0 = \[18] ,
  \[1]  = (f & e) | (~\[8]  | h),
  t2 = ~\[23]  & (~d2 & (~w & ~v)),
  t3 = (~v & u) | ((~v & t) | (~v & s)),
  b0 = \[0] ,
  c0 = \[1] ,
  \[3]  = ~\[8] ,
  d0 = r,
  d2 = \[20]  | ~u,
  \[4]  = (~n & (~j & d)) | ((n & (~j & ~d)) | ((~m & (~j & c)) | ((m & (~j & ~c)) | ((~l & (~j & b)) | ((l & (~j & ~b)) | ((~k & (~j & a)) | (k & (~j & ~a)))))))),
  e0 = \[3] ,
  \[5]  = ~j & ~o,
  f0 = \[4] ,
  \[20]  = ~t | ~s,
  \[6]  = ~j & p,
  g0 = \[5] ,
  \[7]  = ~g | j,
  h0 = \[6] ,
  \[22]  = d2 | ~t3,
  \[8]  = (~t3 & (z & (\x  & w))) | ((z & y) | a0),
  \[10]  = ~q1 & ~s,
  i0 = \[7] ,
  \[23]  = y | \x ,
  \[9]  = ~q & (~h & (f & e)),
  \[11]  = (~q1 & (~\[10]  & ~t)) | (\[10]  & t),
  j0 = \[8] ,
  \[24]  = \[19]  | \x ,
  \[12]  = (~\[20]  & (d2 & ~q1)) | (d2 & (~q1 & u));
endmodule

