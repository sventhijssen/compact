// IWLS benchmark module "count" printed on Wed May 29 16:07:22 2002
module count(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, u, v, w, \x , y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0);
input
  g0,
  h0,
  i0,
  j0,
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  u,
  v,
  w,
  \x ,
  y,
  z,
  a0,
  b0,
  c0,
  d0,
  e0,
  f0;
output
  k0,
  l0,
  m0,
  n0,
  o0,
  p0,
  q0,
  r0,
  s0,
  t0,
  u0,
  v0,
  w0,
  x0,
  y0,
  z0;
wire
  \[26] ,
  \[27] ,
  \[10] ,
  \[11] ,
  \[12] ,
  \[13] ,
  o2,
  \[14] ,
  \[0] ,
  \[15] ,
  \[1] ,
  \[16] ,
  \[2] ,
  \[17] ,
  \[3] ,
  \[18] ,
  \[4] ,
  \[19] ,
  \[5] ,
  \[6] ,
  \[7] ,
  \[8] ,
  y1,
  \[9] ,
  \[20] ,
  \[21] ,
  \[22] ,
  \[23] ,
  e3,
  \[24] ,
  \[25] ;
assign
  \[26]  = \[22]  | e0,
  \[27]  = \[23]  | i0,
  k0 = \[0] ,
  \[10]  = (\[22]  & (e0 & q)) | ((~\[26]  & q) | ((~q & ~f) | s)),
  l0 = \[1] ,
  \[11]  = (\[26]  & (f0 & q)) | ((~e3 & q) | ((~q & ~e) | s)),
  m0 = \[2] ,
  \[12]  = (e3 & (g0 & q)) | ((~\[19]  & q) | ((~q & ~d) | s)),
  n0 = \[3] ,
  \[13]  = (\[19]  & (h0 & q)) | ((~\[23]  & q) | ((~q & ~c) | s)),
  o0 = \[4] ,
  o2 = \[25]  | b0,
  \[14]  = (\[23]  & (i0 & q)) | ((~\[27]  & q) | ((~q & ~b) | s)),
  p0 = \[5] ,
  \[0]  = (u & (r & q)) | ((~\[16]  & q) | ((~q & ~p) | s)),
  \[15]  = (~\[27]  & (~j0 & q)) | ((\[27]  & (j0 & q)) | ((~q & ~a) | s)),
  q0 = \[6] ,
  \[1]  = (\[16]  & (v & q)) | ((~\[20]  & q) | ((~q & ~o) | s)),
  \[16]  = u | r,
  r0 = \[7] ,
  \[2]  = (\[20]  & (w & q)) | ((~\[24]  & q) | ((~q & ~n) | s)),
  \[17]  = y1 | y,
  s0 = \[8] ,
  \[3]  = (\[24]  & (\x  & q)) | ((~y1 & q) | ((~q & ~m) | s)),
  \[18]  = o2 | c0,
  t0 = \[9] ,
  \[4]  = (y1 & (y & q)) | ((~\[17]  & q) | ((~q & ~l) | s)),
  \[19]  = e3 | g0,
  u0 = \[10] ,
  \[5]  = (\[17]  & (z & q)) | ((~\[21]  & q) | ((~q & ~k) | s)),
  v0 = \[11] ,
  \[6]  = (\[21]  & (a0 & q)) | ((~\[25]  & q) | ((~q & ~j) | s)),
  w0 = \[12] ,
  \[7]  = (\[25]  & (b0 & q)) | ((~o2 & q) | ((~q & ~i) | s)),
  x0 = \[13] ,
  \[8]  = (o2 & (c0 & q)) | ((~\[18]  & q) | ((~q & ~h) | s)),
  y0 = \[14] ,
  y1 = \[24]  | \x ,
  \[9]  = (\[18]  & (d0 & q)) | ((~\[22]  & q) | ((~q & ~g) | s)),
  z0 = \[15] ,
  \[20]  = \[16]  | v,
  \[21]  = \[17]  | z,
  \[22]  = \[18]  | d0,
  \[23]  = \[19]  | h0,
  e3 = \[26]  | f0,
  \[24]  = \[20]  | w,
  \[25]  = \[21]  | a0;
endmodule

