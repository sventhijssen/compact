// IWLS benchmark module "cht" printed on Wed May 29 16:07:20 2002
module cht(a, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, \x , y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2, b2, c2, d2, e2, f2);
input
  a,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  t,
  u,
  v,
  w,
  \x ,
  y,
  z,
  a0,
  b0,
  c0,
  d0,
  e0,
  f0,
  g0,
  h0,
  i0,
  j0,
  k0,
  l0,
  m0,
  n0,
  o0,
  p0,
  q0,
  r0,
  s0,
  t0,
  u0,
  v0;
output
  a1,
  a2,
  b1,
  b2,
  c1,
  c2,
  d1,
  d2,
  e1,
  e2,
  f1,
  f2,
  g1,
  h1,
  i1,
  j1,
  k1,
  l1,
  m1,
  n1,
  o1,
  p1,
  q1,
  r1,
  s1,
  t1,
  u1,
  v1,
  w0,
  w1,
  x0,
  x1,
  y0,
  y1,
  z0,
  z1;
wire
  \[5] ,
  \[6] ,
  \[7] ,
  \[8] ,
  \[9] ,
  \[20] ,
  \[21] ,
  \[22] ,
  \[23] ,
  \[24] ,
  \[25] ,
  \[26] ,
  \[27] ,
  \[28] ,
  \[29] ,
  \[30] ,
  \[31] ,
  \[32] ,
  \[33] ,
  \[34] ,
  \[35] ,
  \[36] ,
  \[37] ,
  \[38] ,
  \[39] ,
  \[10] ,
  \[11] ,
  \[12] ,
  \[13] ,
  \[14] ,
  \[15] ,
  \[0] ,
  \[40] ,
  \[16] ,
  \[1] ,
  \[41] ,
  \[17] ,
  \[2] ,
  \[42] ,
  \[18] ,
  \[3] ,
  \[43] ,
  \[19] ,
  \[4] ,
  \[44] ;
assign
  \[5]  = (\[44]  & e) | (\[43]  & r),
  \[6]  = (\[38]  & t) | (\[37]  & s),
  \[7]  = (\[38]  & u) | (\[37]  & t),
  \[8]  = (\[38]  & v) | (\[37]  & u),
  \[9]  = (\[38]  & w) | (\[37]  & v),
  \[20]  = (\[42]  & g0) | (\[40]  & h0),
  \[21]  = (\[42]  & h0) | (\[40]  & i0),
  \[22]  = (\[42]  & i0) | (\[40]  & j0),
  \[23]  = (\[42]  & j0) | (\[40]  & k0),
  \[24]  = (\[42]  & k0) | (\[40]  & l0),
  \[25]  = (\[42]  & l0) | (\[40]  & m0),
  \[26]  = (\[42]  & m0) | (\[40]  & n0),
  \[27]  = (\[40]  & (p & a)) | ((\[42]  & n0) | (\[39]  & o0)),
  \[28]  = (\[41]  & o0) | (\[39]  & p0),
  \[29]  = (\[41]  & p0) | (\[39]  & q0),
  a1 = \[4] ,
  a2 = \[30] ,
  b1 = \[5] ,
  b2 = \[31] ,
  c1 = \[6] ,
  c2 = \[32] ,
  d1 = \[7] ,
  d2 = \[33] ,
  e1 = \[8] ,
  e2 = \[34] ,
  f1 = \[9] ,
  f2 = \[35] ,
  g1 = \[10] ,
  \[30]  = (\[41]  & q0) | (\[39]  & r0),
  h1 = \[11] ,
  \[31]  = (\[41]  & r0) | (\[39]  & s0),
  i1 = \[12] ,
  \[32]  = (\[41]  & s0) | (\[39]  & t0),
  j1 = \[13] ,
  \[33]  = (\[41]  & t0) | (\[39]  & u0),
  k1 = \[14] ,
  \[34]  = (\[41]  & u0) | (\[39]  & v0),
  l1 = \[15] ,
  \[35]  = (\[41]  & v0) | (\[39]  & a),
  m1 = \[16] ,
  \[36]  = p | ~k,
  n1 = \[17] ,
  \[37]  = ~l & ~j,
  o1 = \[18] ,
  \[38]  = ~l & j,
  p1 = \[19] ,
  \[39]  = ~\[36]  & ~l,
  q1 = \[20] ,
  \[10]  = (\[38]  & \x ) | (\[37]  & w),
  r1 = \[21] ,
  \[11]  = (\[38]  & y) | (\[37]  & \x ),
  s1 = \[22] ,
  \[12]  = (\[38]  & z) | (\[37]  & y),
  t1 = \[23] ,
  \[13]  = (\[38]  & a0) | (\[37]  & z),
  u1 = \[24] ,
  \[14]  = (\[38]  & b0) | (\[37]  & a0),
  v1 = \[25] ,
  \[15]  = (\[38]  & c0) | (\[37]  & b0),
  \[0]  = (\[44]  & f) | (\[43]  & m),
  w0 = \[0] ,
  w1 = \[26] ,
  \[40]  = ~l & k,
  \[16]  = (\[38]  & d0) | (\[37]  & c0),
  \[1]  = (\[44]  & g) | (\[43]  & n),
  x0 = \[1] ,
  x1 = \[27] ,
  \[41]  = \[36]  & ~l,
  \[17]  = (\[38]  & e0) | (\[37]  & d0),
  \[2]  = (\[44]  & h) | (\[43]  & o),
  y0 = \[2] ,
  y1 = \[28] ,
  \[42]  = ~l & ~k,
  \[18]  = (\[38]  & f0) | (\[37]  & e0),
  \[3]  = (\[44]  & c) | (\[43]  & p),
  z0 = \[3] ,
  z1 = \[29] ,
  \[43]  = ~l & ~i,
  \[19]  = (\[38]  & a) | (\[37]  & f0),
  \[4]  = (\[44]  & d) | (\[43]  & q),
  \[44]  = ~l & i;
endmodule

