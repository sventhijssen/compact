// IWLS benchmark module "b9" printed on Wed May 29 16:03:33 2002
module b9(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, \x , y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1);
input
  g0,
  h0,
  i0,
  j0,
  k0,
  l0,
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m0,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  t,
  u,
  v,
  w,
  \x ,
  y,
  z,
  n0,
  o0,
  a0,
  b0,
  c0,
  d0,
  e0,
  f0;
output
  g1,
  h1,
  i1,
  j1,
  p0,
  q0,
  r0,
  s0,
  t0,
  u0,
  v0,
  w0,
  x0,
  y0,
  z0,
  a1,
  b1,
  c1,
  d1,
  e1,
  f1;
wire
  f4,
  \[27] ,
  \[28] ,
  j4,
  \[10] ,
  \[11] ,
  \[12] ,
  \[13] ,
  \[0] ,
  \[15] ,
  \[1] ,
  \[16] ,
  \[31] ,
  \[2] ,
  \[17] ,
  \[32] ,
  \[3] ,
  s5,
  \[18] ,
  \[4] ,
  \[34] ,
  \[6] ,
  w2,
  \[7] ,
  \[8] ,
  \[38] ,
  \[9] ,
  \[20] ,
  \[21] ,
  \[23] ,
  \[24] ,
  \[25] ;
assign
  f4 = \[32]  & ~k0,
  g1 = \[17] ,
  h1 = \[18] ,
  \[27]  = ~e0 & ~j,
  i1 = \[11] ,
  \[28]  = ~j0 | ~c0,
  j1 = \[20] ,
  j4 = (c0 & b0) | l0,
  \[10]  = (~\[31]  & (~\[8]  & (h & ~e))) | ((\[34]  & (~\[23]  & f)) | (l0 & (b0 & g))),
  \[11]  = (\[27]  & (\[25]  & (b0 & e))) | ((\[27]  & (\[25]  & c0)) | \[20] ),
  \[12]  = (f4 & (~l0 & (~j0 & ~k))) | ((\[23]  & (~l0 & ~j0)) | ((\[23]  & ~j4) | ((\[23]  & ~b0) | (~b0 & ~k)))),
  \[13]  = ~w2,
  p0 = \[0] ,
  \[0]  = (~\[12]  & ~p) | ~q,
  \[15]  = i0 & (b0 & (a0 & m)),
  q0 = \[1] ,
  \[1]  = ~\[34]  | ~e,
  \[16]  = ~\x  & (w & b),
  r0 = \[2] ,
  \[31]  = f4 | ~b0,
  \[2]  = (~b0 & (~i & e)) | ((\[32]  & e) | ((~d0 & ~c) | ((~i & ~c) | ~\[8] ))),
  \[17]  = ~y & (\x  & (w & b)),
  s0 = \[3] ,
  \[32]  = ~j0 | c0,
  \[3]  = \[38]  | ~v,
  s5 = (~\[28]  & (b0 & (u & (~t & ~s)))) | (l0 & (b0 & (u & (~t & ~s)))),
  \[18]  = ~\[11] ,
  t0 = \[4] ,
  \[4]  = \[38]  | v,
  u0 = j4,
  \[34]  = ~\[31]  | \[24] ,
  v0 = \[6] ,
  \[6]  = ~j4,
  w0 = \[7] ,
  w2 = (~\[24]  & (f4 & (~s5 & c0))) | ((~\[24]  & (~s5 & (~j0 & c0))) | ((~\[24]  & (~s5 & ~b0)) | ((\[23]  & ~s5) | (~s5 & n)))),
  \[7]  = (~h0 & (~f0 & (~z & (~r & (d & a))))) | ((~h0 & (~f0 & (~z & (p & (d & a))))) | ((~m0 & (~h0 & (~f0 & (~r & d)))) | ((~m0 & (~h0 & (~f0 & (p & d)))) | ((~z & (~o & (d & a))) | ((~m0 & (~o & d)) | (z & (~o & d))))))),
  x0 = \[8] ,
  \[8]  = n0 & o0,
  y0 = \[9] ,
  \[38]  = (\[28]  & b0) | ~j4,
  \[9]  = i0 & (b0 & (a0 & l)),
  z0 = \[10] ,
  a1 = \[11] ,
  \[20]  = (\[27]  & (\[21]  & (c0 & ~b0))) | ((\[27]  & (\[25]  & ~j0)) | (\[27]  & (~b0 & ~i))),
  b1 = \[12] ,
  \[21]  = ~\[8]  | ~d0,
  c1 = \[13] ,
  d1 = w2,
  \[23]  = ~\[8]  | e,
  e1 = \[15] ,
  \[24]  = g0 | e0,
  f1 = \[16] ,
  \[25]  = \[21]  | ~i;
endmodule

