// IWLS benchmark module "tcon" printed on Wed May 29 16:09:28 2002
module tcon(a, b, c, d, e, f, g, h, i, k, l, m, n, o, p, q, r, s, t, u, v, w, \x , y, z, a0, b0, c0, d0, e0, f0, g0, h0);
input
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r;
output
  c0,
  d0,
  e0,
  f0,
  g0,
  h0,
  s,
  t,
  u,
  v,
  w,
  \x ,
  y,
  z,
  a0,
  b0;
wire
  \[8] ,
  \[9] ,
  \[10] ,
  \[11] ,
  \[12] ,
  \[13] ,
  \[14] ,
  \[15] ;
assign
  c0 = \[10] ,
  d0 = \[11] ,
  \[8]  = (k & ~i) | (i & a),
  e0 = \[12] ,
  \[9]  = (l & ~i) | (i & b),
  f0 = \[13] ,
  g0 = \[14] ,
  \[10]  = (m & ~i) | (i & c),
  h0 = \[15] ,
  \[11]  = (n & ~i) | (i & d),
  \[12]  = (o & ~i) | (i & e),
  s = k,
  t = l,
  \[13]  = (p & ~i) | (i & f),
  u = m,
  v = n,
  w = o,
  \x  = p,
  y = q,
  z = r,
  \[14]  = (q & ~i) | (i & g),
  \[15]  = (r & ~i) | (i & h),
  a0 = \[8] ,
  b0 = \[9] ;
endmodule

