// IWLS benchmark module "frg2" printed on Wed May 29 16:08:50 2002
module frg2(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, \x , y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2, b2, c2, d2, e2, f2, g2, h2, i2, j2, k2, l2, m2, n2, o2, p2, q2, r2, s2, t2, u2, v2, w2, x2, y2, z2, a3, b3, c3, d3, e3, f3, g3, h3, i3, j3, k3, l3, m3, n3, o3, p3, q3, r3, s3, t3, u3, v3, w3, x3, y3, z3, a4, b4, c4, d4, e4, f4, g4, h4, i4, j4, k4, l4, m4, n4, o4, p4, q4, r4, s4, t4, u4, v4, w4, x4, y4, z4, a5, b5, c5, d5, e5, f5, g5, h5, i5, j5, k5, l5, m5, n5, o5, p5, q5, r5, s5, t5, u5, v5, w5, x5, y5, z5, a6, b6, c6, d6, e6, f6, g6, h6, i6, j6, k6, l6, m6, n6, o6, p6, q6, r6, s6, t6, u6, v6, w6, x6, y6, z6, a7, b7, c7, d7, e7, f7, g7, h7, i7, j7, k7, l7, m7, n7, o7, p7, q7, r7, s7, t7, u7, v7, w7, x7, y7, z7, a8, b8, c8, d8, e8, f8, g8, h8, i8, j8, k8, l8, m8, n8, o8, p8, q8, r8, s8, t8, u8, v8, w8, x8, y8, z8, a9, b9, c9, d9, e9, f9, g9, h9, i9, j9, k9, l9, m9, n9, o9, p9, q9, r9, s9, t9, u9, v9, w9);
input
  z0,
  z1,
  z2,
  z3,
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  t,
  u,
  v,
  w,
  \x ,
  y,
  z,
  a0,
  a1,
  a2,
  a3,
  a4,
  b0,
  b1,
  b2,
  b3,
  b4,
  c0,
  c1,
  c2,
  c3,
  c4,
  d0,
  d1,
  d2,
  d3,
  d4,
  e0,
  e1,
  e2,
  e3,
  e4,
  f0,
  f1,
  f2,
  f3,
  f4,
  g0,
  g1,
  g2,
  g3,
  g4,
  h0,
  h1,
  h2,
  h3,
  h4,
  i0,
  i1,
  i2,
  i3,
  i4,
  j0,
  j1,
  j2,
  j3,
  j4,
  k0,
  k1,
  k2,
  k3,
  k4,
  l0,
  l1,
  l2,
  l3,
  l4,
  m0,
  m1,
  m2,
  m3,
  m4,
  n0,
  n1,
  n2,
  n3,
  n4,
  o0,
  o1,
  o2,
  o3,
  p0,
  p1,
  p2,
  p3,
  q0,
  q1,
  q2,
  q3,
  r1,
  r2,
  r3,
  s0,
  s1,
  s2,
  s3,
  t0,
  t1,
  t2,
  t3,
  u0,
  u1,
  u2,
  u3,
  v0,
  v1,
  v2,
  v3,
  w0,
  w1,
  w2,
  w3,
  x0,
  x1,
  x2,
  x3,
  y0,
  y1,
  y2,
  y3;
output
  z4,
  z5,
  z6,
  z7,
  z8,
  a5,
  a6,
  a7,
  a8,
  a9,
  b5,
  b6,
  b7,
  b8,
  b9,
  c5,
  c6,
  c7,
  c8,
  c9,
  d5,
  d6,
  d7,
  d8,
  d9,
  e5,
  e6,
  e7,
  e8,
  e9,
  f5,
  f6,
  f7,
  f8,
  f9,
  g5,
  g6,
  g7,
  g8,
  g9,
  h5,
  h6,
  h7,
  h8,
  h9,
  i5,
  i6,
  i7,
  i8,
  i9,
  j5,
  j6,
  j7,
  j8,
  j9,
  k5,
  k6,
  k7,
  k8,
  k9,
  l5,
  l6,
  l7,
  l8,
  l9,
  m5,
  m6,
  m7,
  m8,
  m9,
  n5,
  n6,
  n7,
  n8,
  n9,
  o4,
  o5,
  o6,
  o7,
  o8,
  o9,
  p4,
  p5,
  p6,
  p7,
  p8,
  p9,
  q4,
  q5,
  q6,
  q7,
  q8,
  q9,
  r4,
  r5,
  r6,
  r7,
  r8,
  r9,
  s4,
  s5,
  s6,
  s7,
  s8,
  s9,
  t4,
  t5,
  t6,
  t7,
  t8,
  t9,
  u4,
  u5,
  u6,
  u7,
  u8,
  u9,
  v4,
  v5,
  v6,
  v7,
  v8,
  v9,
  w4,
  w5,
  w6,
  w7,
  w8,
  w9,
  x4,
  x5,
  x6,
  x7,
  x8,
  y4,
  y5,
  y6,
  y7,
  y8;
wire
  \[60] ,
  \[145] ,
  \[61] ,
  j25,
  \[146] ,
  j28,
  \[62] ,
  \[63] ,
  \[148] ,
  \[64] ,
  \[149] ,
  r23,
  \[65] ,
  \[66] ,
  \[67] ,
  \[68] ,
  z29,
  \[69] ,
  \[150] ,
  \[0] ,
  \[151] ,
  \[1] ,
  \[152] ,
  \[2] ,
  \[153] ,
  \[3] ,
  c30,
  \[154] ,
  \[4] ,
  \[70] ,
  \[155] ,
  \[71] ,
  \[72] ,
  \[157] ,
  \[7] ,
  \[73] ,
  \[8] ,
  \[74] ,
  \[159] ,
  s23,
  \[9] ,
  \[75] ,
  s28,
  \[76] ,
  \[77] ,
  \[78] ,
  \[79] ,
  \[161] ,
  \[163] ,
  \[164] ,
  \[80] ,
  \[165] ,
  \[81] ,
  l25,
  \[166] ,
  \[82] ,
  \[167] ,
  \[83] ,
  \[168] ,
  t15,
  \[84] ,
  \[169] ,
  t23,
  \[85] ,
  \[86] ,
  \[87] ,
  \[88] ,
  \[89] ,
  \[170] ,
  \[171] ,
  \[10] ,
  \[172] ,
  \[11] ,
  \[173] ,
  \[12] ,
  \[174] ,
  \[13] ,
  \[90] ,
  \[175] ,
  \[14] ,
  \[91] ,
  \[176] ,
  \[15] ,
  \[92] ,
  \[177] ,
  \[16] ,
  \[93] ,
  \[178] ,
  \[17] ,
  \[94] ,
  \[179] ,
  \[18] ,
  \[95] ,
  \[19] ,
  \[96] ,
  \[97] ,
  \[98] ,
  \[100] ,
  \[99] ,
  \[101] ,
  \[102] ,
  \[103] ,
  \[104] ,
  \[181] ,
  \[20] ,
  \[105] ,
  \[21] ,
  \[106] ,
  \[22] ,
  \[107] ,
  \[184] ,
  \[23] ,
  \[108] ,
  \[185] ,
  \[109] ,
  \[186] ,
  \[25] ,
  \[187] ,
  \[26] ,
  \[27] ,
  \[189] ,
  \[28] ,
  \[29] ,
  \[110] ,
  \[111] ,
  \[112] ,
  \[113] ,
  \[114] ,
  \[115] ,
  g25,
  \[116] ,
  \[193] ,
  \[117] ,
  \[118] ,
  \[195] ,
  \[34] ,
  \[119] ,
  \[35] ,
  o29,
  \[36] ,
  \[37] ,
  w16,
  \[38] ,
  \[39] ,
  \[120] ,
  \[121] ,
  \[122] ,
  \[123] ,
  \[124] ,
  \[40] ,
  \[125] ,
  \[41] ,
  \[126] ,
  \[42] ,
  \[127] ,
  \[43] ,
  \[128] ,
  \[44] ,
  \[129] ,
  \[45] ,
  \[46] ,
  \[47] ,
  x15,
  \[48] ,
  \[49] ,
  \[130] ,
  \[131] ,
  a17,
  \[132] ,
  a25,
  \[133] ,
  \[134] ,
  \[135] ,
  \[51] ,
  \[136] ,
  \[52] ,
  \[137] ,
  \[53] ,
  \[138] ,
  \[54] ,
  \[139] ,
  \[55] ,
  \[56] ,
  \[57] ,
  \[58] ,
  \[59] ,
  \[140] ,
  \[141] ,
  \[142] ,
  \[143] ,
  \[144] ;
assign
  \[60]  = (~\[174]  & (~w16 & n1)) | ((~\[174]  & (w16 & o1)) | (~\[189]  & j0)),
  z4 = \[11] ,
  z5 = \[37] ,
  z6 = \[63] ,
  z7 = \[89] ,
  z8 = \[115] ,
  \[145]  = ~\[141]  & \[138] ,
  \[61]  = (~\[174]  & (~w16 & o1)) | ((~\[174]  & (w16 & p1)) | (~\[189]  & i0)),
  j25 = ~\[169]  & ~h4,
  \[146]  = 0,
  j28 = (\[172]  & h1) | ((~s28 & ~h1) | (h1 & ~s0)),
  \[62]  = (~\[174]  & (~w16 & p1)) | ((~\[174]  & (w16 & q1)) | (~\[189]  & h0)),
  \[63]  = (~\[174]  & (~w16 & q1)) | ((~\[174]  & (w16 & r1)) | (~\[189]  & g0)),
  \[148]  = ~z3 | ~y3,
  \[64]  = (~\[174]  & (~w16 & r1)) | ((~\[174]  & (w16 & s1)) | (~\[189]  & f0)),
  \[149]  = ~j1 | z0,
  r23 = ~z29 | m0,
  \[65]  = (~\[174]  & (~w16 & s1)) | ((~\[174]  & (w16 & t1)) | (~\[189]  & e0)),
  \[66]  = (~\[174]  & (~w16 & t1)) | ((~\[174]  & (w16 & u1)) | (~\[189]  & d0)),
  \[67]  = (\[154]  & (~\[139]  & v1)) | ((\[153]  & (~\[139]  & u1)) | ~c30),
  \[68]  = (~\[174]  & (~w16 & v1)) | ((~\[174]  & (w16 & w1)) | (~\[189]  & k0)),
  z29 = ~n0 & t15,
  \[69]  = (~\[174]  & (~w16 & w1)) | ((~\[174]  & (w16 & x1)) | (~\[189]  & l0)),
  \[150]  = ~\[139]  & ~t23,
  \[0]  = ~g1,
  \[151]  = \[139]  | g1,
  \[1]  = (\[185]  & l3) | ((\[152]  & d3) | (~\[22]  & t3)),
  \[152]  = ~s23 & m0,
  \[2]  = (\[185]  & k3) | ((\[152]  & c3) | (~\[21]  & s3)),
  \[153]  = r23 & ~w16,
  \[3]  = (\[185]  & j3) | ((\[152]  & b3) | (~\[20]  & r3)),
  c30 = \[189]  | ~r23,
  \[154]  = r23 & w16,
  \[4]  = (\[185]  & i3) | ((\[152]  & a3) | (~\[19]  & q3)),
  \[70]  = (~\[174]  & (~w16 & x1)) | ((~\[174]  & (w16 & y1)) | (~\[189]  & q)),
  \[155]  = ~h1 | x0,
  \[71]  = (~\[174]  & (~w16 & y1)) | ((~\[174]  & (w16 & z1)) | (~\[189]  & r)),
  \[72]  = (~\[174]  & (~w16 & z1)) | ((~\[174]  & (w16 & a2)) | (~\[189]  & s)),
  \[157]  = ~\[139]  & t23,
  \[7]  = (\[152]  & e3) | (s23 & \[15] ),
  \[73]  = (~\[174]  & (~w16 & a2)) | ((~\[174]  & (w16 & b2)) | (~\[189]  & t)),
  \[8]  = (\[152]  & f3) | (s23 & \[16] ),
  \[74]  = (~\[174]  & (~w16 & b2)) | ((~\[174]  & (w16 & c2)) | (~\[189]  & u)),
  \[159]  = a4 | ~z3,
  s23 = (~l0 & k0) | (l0 & ~k0),
  \[9]  = (\[152]  & g3) | (s23 & \[17] ),
  \[75]  = (~\[174]  & (~w16 & c2)) | ((~\[174]  & (w16 & d2)) | (~\[189]  & v)),
  s28 = (l1 & (~k1 & (~j1 & (~i1 & w0)))) | ((~\[179]  & (~l1 & (k1 & ~i1))) | ((~\[173]  & (j1 & (~i1 & u0))) | (~g25 & (i1 & t0)))),
  \[76]  = (~\[174]  & (~w16 & d2)) | ((~\[174]  & (w16 & e2)) | (~\[189]  & w)),
  \[77]  = (~\[174]  & (~w16 & e2)) | ((~\[174]  & (w16 & f2)) | (~\[189]  & \x )),
  \[78]  = (~\[174]  & (~w16 & f2)) | ((~\[174]  & (w16 & g2)) | (~\[189]  & y)),
  \[79]  = (~\[174]  & (~w16 & g2)) | ((~\[174]  & (w16 & h2)) | (~\[189]  & z)),
  \[161]  = \[148]  | (b4 | a4),
  \[163]  = \[150]  & ~w16,
  \[164]  = ~r23 & (s23 & k0),
  \[80]  = (~\[174]  & (~w16 & h2)) | ((~\[174]  & (w16 & i2)) | (~\[189]  & a0)),
  \[165]  = g4 | ~f4,
  \[81]  = (~\[174]  & (~w16 & i2)) | ((~\[174]  & (w16 & j2)) | (~\[189]  & b0)),
  l25 = (l1 & ~b1) | (~\[176]  | (~\[175]  | (~\[155]  | ~\[149] ))),
  \[166]  = \[161]  | c4,
  \[82]  = (~\[174]  & (~w16 & j2)) | ((~\[174]  & (w16 & k2)) | (~\[189]  & c0)),
  \[167]  = \[150]  & w16,
  \[83]  = (\[164]  & (~\[139]  & i)) | ((\[154]  & (~\[139]  & l2)) | ((\[153]  & (~\[139]  & k2)) | (\[142]  & (~\[139]  & a)))),
  \[168]  = ~j25 & n4,
  t15 = ~\[172]  & ~h1,
  \[84]  = (\[164]  & (~\[139]  & j)) | ((\[154]  & (~\[139]  & m2)) | ((\[153]  & (~\[139]  & l2)) | (\[142]  & (~\[139]  & b)))),
  \[169]  = \[165]  | ~e4,
  t23 = ~r23 & ~s23,
  \[85]  = (\[164]  & (~\[139]  & k)) | ((\[154]  & (~\[139]  & n2)) | ((\[153]  & (~\[139]  & m2)) | (\[142]  & (~\[139]  & c)))),
  \[86]  = (\[164]  & (~\[139]  & l)) | ((\[154]  & (~\[139]  & o2)) | ((\[153]  & (~\[139]  & n2)) | (\[142]  & (~\[139]  & d)))),
  \[87]  = (\[164]  & (~\[139]  & m)) | ((\[154]  & (~\[139]  & p2)) | ((\[153]  & (~\[139]  & o2)) | (\[142]  & (~\[139]  & e)))),
  \[88]  = (\[164]  & (~\[139]  & n)) | ((\[154]  & (~\[139]  & q2)) | ((\[153]  & (~\[139]  & p2)) | (\[142]  & (~\[139]  & f)))),
  \[89]  = (\[164]  & (~\[139]  & o)) | ((\[154]  & (~\[139]  & r2)) | ((\[153]  & (~\[139]  & q2)) | (\[142]  & (~\[139]  & g)))),
  \[170]  = k4 | n0,
  \[171]  = k4 | ~m1,
  \[10]  = (\[152]  & h3) | (s23 & \[18] ),
  \[172]  = g25 | i1,
  \[11]  = (\[152]  & i3) | (s23 & \[19] ),
  \[173]  = l1 | k1,
  \[12]  = (\[152]  & j3) | (s23 & \[20] ),
  \[174]  = \[139]  | z29,
  \[13]  = (\[152]  & k3) | (s23 & \[21] ),
  \[90]  = (\[164]  & (~\[139]  & p)) | ((\[154]  & (~\[139]  & s2)) | ((\[153]  & (~\[139]  & r2)) | (\[142]  & (~\[139]  & h)))),
  \[175]  = ~k1 | a1,
  \[14]  = (\[152]  & l3) | (s23 & \[22] ),
  \[91]  = (\[167]  & t2) | ((\[163]  & s2) | (\[157]  & i)),
  \[176]  = ~i1 | y0,
  \[15]  = m0 & m3,
  \[92]  = (\[167]  & u2) | ((\[163]  & t2) | (\[157]  & j)),
  \[177]  = ~l25 | ~k4,
  \[16]  = m0 & n3,
  \[93]  = (\[167]  & v2) | ((\[163]  & u2) | (\[157]  & k)),
  \[178]  = j25 | d4,
  \[17]  = m0 & o3,
  \[94]  = (\[167]  & w2) | ((\[163]  & v2) | (\[157]  & l)),
  \[179]  = j1 | ~v0,
  \[18]  = m0 & p3,
  \[95]  = (\[167]  & x2) | ((\[163]  & w2) | (\[157]  & m)),
  \[19]  = m0 & q3,
  \[96]  = (\[167]  & y2) | ((\[163]  & x2) | (\[157]  & n)),
  \[97]  = (\[167]  & z2) | ((\[163]  & y2) | (\[157]  & o)),
  \[98]  = (\[163]  & z2) | (\[157]  & p),
  \[100]  = (\[145]  & c3) | (\[143]  & b3),
  \[99]  = (\[145]  & b3) | (\[143]  & a3),
  \[101]  = (\[145]  & d3) | (\[143]  & c3),
  \[102]  = (\[145]  & e3) | (\[143]  & d3),
  \[103]  = (\[145]  & f3) | (\[143]  & e3),
  \[104]  = (\[145]  & g3) | (\[143]  & f3),
  \[181]  = \[151]  | z29,
  \[20]  = m0 & r3,
  \[105]  = (\[145]  & h3) | (\[143]  & g3),
  \[21]  = m0 & s3,
  \[106]  = (\[145]  & i3) | (\[143]  & h3),
  \[22]  = m0 & t3,
  \[107]  = (\[145]  & j3) | (\[143]  & i3),
  \[184]  = ~\[139]  & ~x15,
  \[23]  = ~j4 & g1,
  \[108]  = (\[145]  & k3) | (\[143]  & j3),
  \[185]  = s23 & m0,
  \[109]  = (\[145]  & l3) | (\[143]  & k3),
  \[186]  = ~\[151] ,
  \[25]  = \[170]  | ~h1,
  \[187]  = \[129]  | ~e4,
  \[26]  = \[170]  | ~i1,
  \[27]  = \[170]  | ~j1,
  \[189]  = \[139]  | ~z29,
  \[28]  = \[170]  | ~k1,
  \[29]  = \[170]  | ~l1,
  \[110]  = (\[145]  & m3) | (\[143]  & l3),
  \[111]  = (\[145]  & n3) | (\[143]  & m3),
  \[112]  = (\[145]  & o3) | (\[143]  & n3),
  \[113]  = (\[145]  & p3) | (\[143]  & o3),
  \[114]  = (\[145]  & q3) | (\[143]  & p3),
  \[115]  = (\[145]  & r3) | (\[143]  & q3),
  g25 = \[173]  | j1,
  \[116]  = (\[145]  & s3) | (\[143]  & r3),
  \[193]  = \[178]  | ~\[128] ,
  \[117]  = (\[145]  & t3) | (\[143]  & s3),
  \[118]  = (\[145]  & u3) | (\[143]  & t3),
  \[195]  = ~\[139]  & m1,
  \[34]  = (~\[166]  & \[51] ) | (\[166]  & n1),
  \[119]  = (\[145]  & v3) | (\[143]  & u3),
  \[35]  = \[171]  | ~h1,
  o29 = ~a17 & (~x3 & y3),
  \[36]  = \[171]  | ~i1,
  \[37]  = \[171]  | ~j1,
  w16 = ~a17 & l4,
  \[38]  = \[171]  | ~k1,
  \[39]  = \[171]  | ~l1,
  \[120]  = (\[145]  & w3) | (\[143]  & v3),
  \[121]  = (~j25 & (~j28 & \[138] )) | (\[143]  & w3),
  \[122]  = (~\[174]  & (~w16 & x3)) | (~\[174]  & (w16 & ~x3)),
  \[123]  = (~o29 & (w16 & \[122] )) | ((~o29 & y3) | ((o29 & ~w16) | \[174] )),
  \[124]  = (\[148]  & (o29 & ~\[123] )) | ((~\[148]  & ~w16) | ((~o29 & z3) | \[174] )),
  \[40]  = ~l4 | ~h1,
  \[125]  = (~\[159]  & (\[154]  & (~\[139]  & o29))) | ((\[148]  & (~\[139]  & (r23 & a4))) | ((~\[139]  & (~o29 & (r23 & a4))) | ((\[153]  & (~\[139]  & a4)) | (\[157]  | ~c30)))),
  \[41]  = ~l4 | ~i1,
  \[126]  = (~\[174]  & (\[124]  & b4)) | ((\[159]  & (~\[124]  & b4)) | ((~\[161]  & ~\[124] ) | ~c30)),
  \[42]  = ~l4 | ~j1,
  \[127]  = (~\[139]  & (c30 & (\[124]  & c4))) | ((\[159]  & (~\[124]  & c4)) | ((~\[124]  & (c4 & b4)) | (~\[139]  & ~r23))),
  \[43]  = ~l4 | ~k1,
  \[128]  = (~\[178]  & (\[138]  & ~g1)) | ((\[177]  & (~\[151]  & d4)) | ((~\[151]  & (j25 & d4)) | ~\[189] )),
  \[44]  = ~l4 | ~l1,
  \[129]  = (~\[193]  & ~e4) | ((\[193]  & e4) | \[181] ),
  \[45]  = ~h1,
  \[46]  = ~i1,
  \[47]  = ~j1,
  x15 = ~z29 | e1,
  a5 = \[12] ,
  a6 = \[38] ,
  a7 = \[64] ,
  a8 = \[90] ,
  a9 = \[116] ,
  \[48]  = ~k1,
  b5 = \[13] ,
  b6 = \[39] ,
  b7 = \[65] ,
  b8 = \[91] ,
  b9 = \[117] ,
  \[49]  = ~l1,
  c5 = \[14] ,
  c6 = \[40] ,
  c7 = \[66] ,
  c8 = \[92] ,
  c9 = \[118] ,
  d5 = \[15] ,
  d6 = \[41] ,
  d7 = \[67] ,
  d8 = \[93] ,
  d9 = \[119] ,
  e5 = \[16] ,
  e6 = \[42] ,
  e7 = \[68] ,
  e8 = \[94] ,
  e9 = \[120] ,
  \[130]  = (~\[187]  & ~f4) | ((\[187]  & f4) | \[181] ),
  f5 = \[17] ,
  f6 = \[43] ,
  f7 = \[69] ,
  f8 = \[95] ,
  f9 = \[121] ,
  \[131]  = (~\[181]  & (\[130]  & g4)) | ((~\[181]  & (g4 & ~f4)) | ((\[181]  & (~s23 & \[128] )) | ((~\[165]  & ~\[130] ) | (~r23 & \[128] )))),
  g5 = \[18] ,
  g6 = \[44] ,
  g7 = \[70] ,
  g8 = \[96] ,
  g9 = \[122] ,
  a17 = ~\[166]  & ~x3,
  \[132]  = (~\[181]  & (\[169]  & h4)) | ((~\[181]  & (~\[138]  & h4)) | ((~\[181]  & (~\[128]  & h4)) | ~c30)),
  h5 = \[19] ,
  h6 = \[45] ,
  h7 = \[71] ,
  h8 = \[97] ,
  h9 = \[123] ,
  a25 = \[139]  | ~l25,
  \[133]  = (~\[139]  & (w16 & (~i4 & n1))) | (~\[139]  & (w16 & (i4 & ~n1))),
  i5 = \[20] ,
  i6 = \[46] ,
  i7 = \[72] ,
  i8 = \[98] ,
  i9 = \[124] ,
  \[134]  = (\[168]  & (~\[151]  & (\[145]  & (~j28 & ~j4)))) | ((~\[151]  & (~\[145]  & j4)) | ((~\[151]  & (j28 & j4)) | (~\[151]  & (~n4 & j4)))),
  j5 = \[21] ,
  j6 = \[47] ,
  j7 = \[73] ,
  j8 = \[99] ,
  j9 = \[125] ,
  \[135]  = \[195]  & ~\[166] ,
  \[51]  = (~i4 & ~f1) | (i4 & f1),
  k5 = \[22] ,
  k6 = \[48] ,
  k7 = \[74] ,
  k8 = \[100] ,
  k9 = \[126] ,
  \[136]  = \[195]  & ~a17,
  \[52]  = ~\[166]  & x3,
  l5 = \[23] ,
  l6 = \[49] ,
  l7 = \[75] ,
  l8 = \[101] ,
  l9 = \[127] ,
  \[137]  = (\[168]  & \[53] ) | (l25 & \[53] ),
  \[53]  = (\[168]  & (~\[139]  & ~l25)) | (~\[151]  & (j25 & d4)),
  m5 = m4,
  m6 = k4,
  m7 = \[76] ,
  m8 = \[102] ,
  m9 = \[128] ,
  \[138]  = ~a25 & k4,
  \[54]  = (\[186]  & h1) | (\[184]  & ~\[144] ),
  n5 = \[25] ,
  n6 = \[51] ,
  n7 = \[77] ,
  n8 = \[103] ,
  n9 = \[129] ,
  \[139]  = q0 | ~o0,
  \[55]  = (\[184]  & (~d1 & c1)) | (\[186]  & i1),
  o4 = \[0] ,
  o5 = \[26] ,
  o6 = \[52] ,
  o7 = \[78] ,
  o8 = \[104] ,
  o9 = \[130] ,
  \[56]  = (\[184]  & (d1 & ~c1)) | (\[186]  & j1),
  p4 = \[1] ,
  p5 = \[27] ,
  p6 = \[53] ,
  p7 = \[79] ,
  p8 = \[105] ,
  p9 = \[131] ,
  \[57]  = (\[184]  & (d1 & c1)) | (\[186]  & k1),
  q4 = \[2] ,
  q5 = \[28] ,
  q6 = \[54] ,
  q7 = \[80] ,
  q8 = \[106] ,
  q9 = \[132] ,
  \[58]  = (~\[189]  & (~\[144]  & x15)) | (~\[151]  & l1),
  r4 = \[3] ,
  r5 = \[29] ,
  r6 = \[55] ,
  r7 = \[81] ,
  r8 = \[107] ,
  r9 = \[133] ,
  \[59]  = (~\[139]  & (~m1 & (p0 & ~n0))) | (\[195]  & ~\[53] ),
  s4 = \[4] ,
  s5 = \[34] ,
  s6 = \[56] ,
  s7 = \[82] ,
  s8 = \[108] ,
  s9 = \[134] ,
  t4 = u3,
  t5 = \[34] ,
  t6 = \[57] ,
  t7 = \[83] ,
  t8 = \[109] ,
  t9 = \[135] ,
  u4 = v3,
  u5 = \[34] ,
  u6 = \[58] ,
  u7 = \[84] ,
  u8 = \[110] ,
  u9 = \[136] ,
  \[140]  = 0,
  v4 = \[7] ,
  v5 = \[34] ,
  v6 = \[59] ,
  v7 = \[85] ,
  v8 = \[111] ,
  v9 = \[137] ,
  \[141]  = (\[173]  & j1) | ((\[172]  & h1) | ((g25 & i1) | ((l1 & k1) | (j25 | t15)))),
  w4 = \[8] ,
  w5 = \[34] ,
  w6 = \[60] ,
  w7 = \[86] ,
  w8 = \[112] ,
  w9 = \[138] ,
  \[142]  = (~r23 & l0) | t23,
  x4 = \[9] ,
  x5 = \[35] ,
  x6 = \[61] ,
  x7 = \[87] ,
  x8 = \[113] ,
  \[143]  = (\[177]  & ~\[139] ) | (\[141]  & ~\[139] ),
  y4 = \[10] ,
  y5 = \[36] ,
  y6 = \[62] ,
  y7 = \[88] ,
  y8 = \[114] ,
  \[144]  = d1 | c1;
endmodule

