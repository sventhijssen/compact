// IWLS benchmark module "b9" printed on Wed May 29 16:03:33 2002
module b9(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, \x , y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1);
input
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  t,
  u,
  v,
  w,
  \x ,
  y,
  z,
  a0,
  b0,
  c0,
  d0,
  e0,
  f0,
  g0,
  h0,
  i0,
  j0,
  k0,
  l0,
  m0,
  n0,
  o0;
output
  a1,
  b1,
  c1,
  d1,
  e1,
  f1,
  g1,
  h1,
  i1,
  j1,
  p0,
  q0,
  r0,
  s0,
  t0,
  u0,
  v0,
  w0,
  x0,
  y0,
  z0;
wire
  \[6] ,
  \[7] ,
  \[8] ,
  \[9] ,
  \[20] ,
  a5,
  b5,
  c5,
  d4,
  d5,
  e4,
  e5,
  f3,
  f4,
  g2,
  g3,
  g5,
  h2,
  h4,
  i2,
  i3,
  i4,
  i5,
  j3,
  j4,
  j5,
  k2,
  k3,
  l2,
  l4,
  m2,
  m3,
  m4,
  m5,
  n3,
  n5,
  o3,
  o5,
  p5,
  q2,
  \[10] ,
  q3,
  q5,
  r2,
  \[11] ,
  r4,
  r5,
  s2,
  \[12] ,
  s3,
  s4,
  s5,
  t2,
  \[13] ,
  t3,
  t4,
  t5,
  u2,
  u4,
  u5,
  v2,
  \[15] ,
  v4,
  v5,
  \[0] ,
  w2,
  \[16] ,
  w3,
  w5,
  \[1] ,
  x2,
  \[17] ,
  x3,
  x4,
  \[2] ,
  \[18] ,
  y3,
  \[3] ,
  z3,
  \[4] ;
assign
  \[6]  = ~j4,
  \[7]  = (~m0 & ~u2) | (~v2 & ~u2),
  \[8]  = ~a5,
  \[9]  = ~x2,
  \[20]  = (~t2 & ~s2) | (~n0 & ~s2),
  a1 = \[11] ,
  a5 = ~n0 | ~o0,
  b1 = \[12] ,
  b5 = g0 | e0,
  c1 = \[13] ,
  c5 = ~o0 | e,
  d1 = w2,
  d4 = \x  | (~w | ~b),
  d5 = (~t5 & ~b5) | (~b0 & ~b5),
  e1 = \[15] ,
  e4 = y | (~\x  | (~w | ~b)),
  e5 = ~d5 & (~c5 & ~n),
  f1 = \[16] ,
  f3 = ~k3 & v,
  f4 = (~k0 & ~j0) | (~k0 & c0),
  g1 = \[17] ,
  g2 = ~m2 | (~l2 | ~k2),
  g3 = ~k3 & ~v,
  g5 = ~j0 | c0,
  h1 = \[18] ,
  h2 = ~i2 & o0,
  h4 = f4 | (~b0 | (~h | e)),
  i1 = \[11] ,
  i2 = ~d0 | ~i,
  i3 = w5 | (~b0 | ~m),
  i4 = ~f4 & o0,
  i5 = ~l0 | (~g | ~b0),
  j1 = \[20] ,
  j3 = j0 & c0,
  j4 = (c0 & b0) | l0,
  j5 = ~m5 | (~n0 | (~f | e)),
  k2 = ~e0 & ~j,
  k3 = (~j3 & ~l0) | ((~j3 & b0) | (~l0 & ~b0)),
  l2 = ~j0 | (c0 | (~b0 | e)),
  l4 = r & ~p,
  m2 = ~n3 | b0,
  m3 = (~v5 & e) | ~q3,
  m4 = ~h0 & (~f0 & ~l4),
  m5 = ~p5 | ~o5,
  n3 = j0 & (~c0 & i),
  n5 = (~n0 & ~h4) | (~o0 & ~h4),
  o3 = ~d0 | ~i,
  o5 = ~b0 | ~i4,
  p0 = \[0] ,
  p5 = ~o0 | ~q5,
  q0 = \[1] ,
  q2 = j0 & c0,
  \[10]  = n5 | (~j5 | ~i5),
  q3 = ~o3 | c,
  q5 = g0 | e0,
  r0 = \[2] ,
  r2 = ~q2 & ~l0,
  \[11]  = (~h2 & ~g2) | (~n0 & ~g2),
  r4 = ~u | (t | s),
  r5 = (~j0 & ~l0) | (~c0 & ~l0),
  s0 = \[3] ,
  s2 = ~s3 | (~t3 | (e0 | j)),
  \[12]  = (~n0 & ~u5) | (~t4 & ~u5),
  s3 = ~j0 | (c0 | ~i),
  s4 = (~v4 & ~x4) | (~b0 & ~x4),
  s5 = ~r5 & (~r4 & b0),
  t0 = \[4] ,
  t2 = o0 & (d0 & i),
  \[13]  = ~w2,
  t3 = ~b0 | ~j0,
  t4 = ~s4 & o0,
  t5 = (k0 & j0) | ~c0,
  u0 = j4,
  u2 = (~m4 & o) | ~d,
  u4 = (~k0 & ~j0) | (~k0 & c0),
  u5 = ~r2 & b0,
  v0 = \[6] ,
  v2 = (~z & ~a) | ((z & o) | (o & ~a)),
  \[15]  = ~i3,
  v4 = ~e & ~u4,
  v5 = (~g5 & b0) | (~g5 & i),
  \[0]  = (~\[12]  & ~p) | ~q,
  w0 = \[7] ,
  w2 = (~e5 & ~s5) | (~n0 & ~s5),
  \[16]  = ~d4,
  w3 = ~k0 | (~b0 | ~e),
  w5 = ~a0 | ~i0,
  \[1]  = ~z3,
  x0 = \[8] ,
  x2 = w5 | (~b0 | ~l),
  \[17]  = ~e4,
  x3 = ~j0 | (c0 | (~b0 | ~e)),
  x4 = k & ~e,
  \[2]  = m3 | (~o0 | ~n0),
  y0 = \[9] ,
  \[18]  = ~\[11] ,
  y3 = (~g0 & ~e0) | ~e,
  \[3]  = ~f3,
  z0 = \[10] ,
  z3 = ~y3 | (~x3 | ~w3),
  \[4]  = ~g3;
endmodule

