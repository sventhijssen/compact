// IWLS benchmark module "ldd" printed on Wed May 29 16:09:11 2002
module ldd(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, \x , y, z, a0, b0);
input
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i;
output
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  t,
  u,
  v,
  w,
  \x ,
  y,
  z,
  a0,
  b0;
wire
  \[13] ,
  \[14] ,
  \[15] ,
  \[16] ,
  o1,
  \[17] ,
  p1,
  \[18] ,
  q1,
  r1,
  s1,
  \[0] ,
  t1,
  \[1] ,
  u1,
  \[2] ,
  v1,
  \[3] ,
  w1,
  \[4] ,
  x1,
  \[5] ,
  y1,
  \[6] ,
  z1,
  \[7] ,
  \[8] ,
  \[10] ,
  \[9] ,
  \[11] ,
  \[12] ;
assign
  \[13]  = \[11]  | (\[10]  | (\[9]  | (\[8]  | (s1 | (r1 | (q1 | p1)))))),
  \[14]  = \[11]  | (\[10]  | (\[9]  | (\[8]  | (s1 | (r1 | (q1 | p1)))))),
  \[15]  = \[10]  | (\[8]  | (s1 | q1)),
  \[16]  = \[11]  | (\[8]  | (s1 | p1)),
  o1 = ~i & (~c & (~b & a)),
  \[17]  = \[11]  | (s1 | (r1 | q1)),
  p1 = h & (~g & (~f & (~e & (~d & (~c & (~b & ~a)))))),
  \[18]  = d & (~c & (~b & ~a)),
  q1 = g & (~f & (~e & (~d & (~c & (~b & ~a))))),
  j = \[0] ,
  k = \[1] ,
  l = \[2] ,
  m = \[3] ,
  n = \[4] ,
  o = \[5] ,
  p = \[6] ,
  q = \[7] ,
  r = \[8] ,
  s = \[9] ,
  r1 = f & (~e & (~d & (~c & (~b & ~a)))),
  t = \[10] ,
  u = \[11] ,
  v = \[12] ,
  w = \[13] ,
  \x  = \[14] ,
  y = \[15] ,
  z = \[16] ,
  s1 = e & (~d & (~c & (~b & ~a))),
  \[0]  = w1 | (v1 | (\[11]  | (z1 | (\[10]  | (o1 | (\[9]  | (\[8]  | (u1 | (q1 | p1))))))))),
  a0 = \[17] ,
  t1 = ~i & (c & (~b & ~a)),
  \[1]  = w1 | (v1 | (\[11]  | (\[10]  | (\[9]  | (y1 | (\[8]  | (x1 | (u1 | (s1 | r1))))))))),
  b0 = \[18] ,
  u1 = i & (c & (~b & ~a)),
  \[2]  = w1 | (z1 | (\[10]  | (\[9]  | (y1 | (\[8]  | (u1 | (t1 | (\[18]  | (r1 | p1))))))))),
  v1 = ~i & (~c & (b & a)),
  \[3]  = \[11]  | (z1 | (\[9]  | (y1 | (\[8]  | x1)))),
  w1 = i & (~c & (b & a)),
  \[4]  = \[10]  | o1,
  x1 = ~i & (~c & (b & ~a)),
  \[5]  = w1 | v1,
  y1 = ~i & (c & (b & ~a)),
  \[6]  = u1 | t1,
  z1 = ~i & (c & (~b & a)),
  \[7]  = (~h & (~g & (~f & (~e & (~d & (~c & (~b & ~a))))))) | (\[18]  | (s1 | (r1 | (q1 | p1)))),
  \[8]  = i & (~c & (b & ~a)),
  \[10]  = i & (~c & (~b & a)),
  \[9]  = i & (c & (b & ~a)),
  \[11]  = i & (c & (~b & a)),
  \[12]  = \[11]  | (z1 | (\[10]  | (\[9]  | (\[8]  | (s1 | (r1 | (q1 | p1)))))));
endmodule

