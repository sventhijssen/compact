// IWLS benchmark module "sct" printed on Wed May 29 16:09:28 2002
module sct(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, \x , y, z, a0, b0, c0, d0, e0, f0, g0, h0);
input
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s;
output
  t,
  u,
  v,
  w,
  \x ,
  y,
  z,
  a0,
  b0,
  c0,
  d0,
  e0,
  f0,
  g0,
  h0;
wire
  \[14] ,
  \[15] ,
  \[16] ,
  \[17] ,
  \[18] ,
  \[0] ,
  \[1] ,
  \[2] ,
  \[3] ,
  \[4] ,
  \[5] ,
  \[20] ,
  \[6] ,
  \[21] ,
  \[7] ,
  \[22] ,
  \[8] ,
  \[10] ,
  \[23] ,
  \[9] ,
  \[12] ;
assign
  \[14]  = e & r,
  \[15]  = \[16]  & e,
  \[16]  = ~\[12]  | ~q,
  \[17]  = ~\[15] ,
  \[18]  = ~\[5]  | j,
  t = \[0] ,
  u = \[1] ,
  v = \[2] ,
  w = \[3] ,
  \x  = \[4] ,
  y = \[5] ,
  z = \[6] ,
  \[0]  = (~o & ~b) | (~c & b),
  a0 = \[7] ,
  \[1]  = (~s & ~f) | ((p & ~f) | (f & ~e)),
  b0 = \[8] ,
  \[2]  = ~\[17]  & ~g,
  c0 = \[9] ,
  \[3]  = (\[16]  & (~\[2]  & (~h & e))) | (\[2]  & h),
  d0 = \[10] ,
  \[4]  = (\[15]  & (~\[3]  & (~i & h))) | ((\[3]  & i) | (\[2]  & i)),
  e0 = c,
  \[5]  = (~\[20]  & ~j) | ((\[20]  & j) | \[17] ),
  f0 = \[12] ,
  \[20]  = \[4]  | ~i,
  \[6]  = (~\[18]  & ~k) | ((\[18]  & k) | \[17] ),
  g0 = e,
  \[21]  = ~\[6]  | k,
  \[7]  = (~\[21]  & ~l) | ((\[21]  & l) | \[17] ),
  h0 = \[14] ,
  \[22]  = ~\[7]  | l,
  \[8]  = (~\[22]  & ~m) | ((\[22]  & m) | \[17] ),
  \[10]  = (~\[18]  & (\[15]  & (~n & (~m & (~l & ~k))))) | ((~\[18]  & (\[15]  & a)) | (~\[16]  & o)),
  \[23]  = ~\[8]  | m,
  \[9]  = (~\[23]  & ~n) | ((\[23]  & n) | \[17] ),
  \[12]  = (q & (e & ~c)) | (d & e);
endmodule

