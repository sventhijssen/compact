// IWLS benchmark module "c8" printed on Wed May 29 16:07:19 2002
module c8(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, u, v, w, \x , y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0);
input
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  u,
  v,
  w,
  \x ,
  y,
  z,
  a0,
  b0,
  c0;
output
  g0,
  h0,
  i0,
  j0,
  k0,
  l0,
  m0,
  n0,
  o0,
  p0,
  q0,
  r0,
  s0,
  t0,
  u0,
  d0,
  e0,
  f0;
wire
  g2,
  h2,
  i2,
  j2,
  k2,
  \[10] ,
  \[11] ,
  m2,
  \[12] ,
  n2,
  \[13] ,
  o2,
  \[14] ,
  p2,
  \[0] ,
  \[15] ,
  q2,
  \[1] ,
  \[16] ,
  \[2] ,
  \[17] ,
  s2,
  \[3] ,
  t2,
  \[4] ,
  u1,
  u2,
  \[5] ,
  v1,
  v2,
  \[6] ,
  w1,
  w2,
  \[7] ,
  y1,
  y2,
  \[9] ,
  z1,
  z2,
  a2,
  a3,
  b3,
  c2,
  c3,
  d2,
  d3,
  e2;
assign
  g0 = \[3] ,
  g2 = ~i2 | (r | (u | v)),
  h0 = \[4] ,
  h2 = (~s & (~q & ~m)) | ((s & (~q & ~e)) | (~q & (~m & ~e))),
  i0 = \[5] ,
  i2 = ~w & ~\x ,
  j0 = \[6] ,
  j2 = ~u & ~v,
  k0 = \[7] ,
  k2 = ~w & (~\x  & (~y & z)),
  \[10]  = (~v1 & ~u1) | ((~v1 & ~q) | (~v1 & v)),
  l0 = c0,
  \[11]  = (~z1 & (~y1 & ~w1)) | ((~z1 & (~y1 & r)) | ((~z1 & (~y1 & u)) | ((~z1 & (w & ~w1)) | ((~z1 & (w & r)) | ((~z1 & (w & u)) | (~z1 & ~q)))))),
  m0 = \[9] ,
  m2 = ~o2 | (r | (u | v)),
  \[12]  = (~d2 & (~c2 & ~a2)) | ((~d2 & (~c2 & r)) | ((~d2 & (~c2 & u)) | ((~d2 & (\x  & ~a2)) | ((~d2 & (\x  & r)) | ((~d2 & (\x  & u)) | (~d2 & ~q)))))),
  n0 = \[10] ,
  n2 = (~s & (~q & ~n)) | ((s & (~q & ~f)) | (~q & (~n & ~f))),
  \[13]  = (~h2 & (~g2 & ~e2)) | ((~h2 & (~g2 & r)) | ((~h2 & (~g2 & u)) | ((~h2 & (y & ~e2)) | ((~h2 & (y & r)) | ((~h2 & (y & u)) | (~h2 & ~q)))))),
  o0 = \[11] ,
  o2 = ~w & (~\x  & ~y),
  \[14]  = (~n2 & (~m2 & ~k2)) | ((~n2 & (~m2 & ~j2)) | ((~n2 & (~m2 & r)) | ((~n2 & (z & ~k2)) | ((~n2 & (z & ~j2)) | ((~n2 & (z & r)) | (~n2 & ~q)))))),
  p0 = \[12] ,
  p2 = ~u & (~v & ~w),
  \[0]  = (~c0 & ~u) | ((c0 & ~i) | (~u & ~i)),
  \[15]  = (~t2 & (~s2 & ~q2)) | ((~t2 & (~s2 & ~p2)) | ((~t2 & (~s2 & r)) | ((~t2 & (a0 & ~q2)) | ((~t2 & (a0 & ~p2)) | ((~t2 & (a0 & r)) | (~t2 & ~q)))))),
  q0 = \[13] ,
  q2 = ~\x  & (~y & (~z & a0)),
  \[1]  = (~c0 & ~v) | ((c0 & ~j) | (~v & ~j)),
  \[16]  = (~z2 & (~y2 & ~w2)) | ((~z2 & (~y2 & ~v2)) | ((~z2 & (~y2 & r)) | ((~z2 & (b0 & ~w2)) | ((~z2 & (b0 & ~v2)) | ((~z2 & (b0 & r)) | (~z2 & ~q)))))),
  r0 = \[14] ,
  \[2]  = (~c0 & ~w) | ((c0 & ~k) | (~w & ~k)),
  \[17]  = (~d3 & (~c3 & (~r & q))) | (c0 & (r & q)),
  s0 = \[15] ,
  s2 = ~u2 | (r | (u | v)),
  \[3]  = (~c0 & ~\x ) | ((c0 & ~l) | (~\x  & ~l)),
  t0 = \[16] ,
  t2 = (~s & (~q & ~o)) | ((s & (~q & ~g)) | (~q & (~o & ~g))),
  \[4]  = (~c0 & ~y) | ((c0 & ~m) | (~y & ~m)),
  u0 = \[17] ,
  u1 = r | u,
  u2 = ~w & (~\x  & (~y & ~z)),
  \[5]  = (~c0 & ~z) | ((c0 & ~n) | (~z & ~n)),
  v1 = (v & (~u & (~r & q))) | ((~s & (~q & ~j)) | (s & (~q & ~b))),
  v2 = ~u & (~v & (~w & ~\x )),
  \[6]  = (~c0 & ~a0) | ((c0 & ~o) | (~a0 & ~o)),
  w1 = ~v & w,
  w2 = ~y & (~z & (~a0 & b0)),
  \[7]  = (~c0 & ~b0) | ((c0 & ~p) | (~b0 & ~p)),
  y1 = r | (u | v),
  y2 = ~b3 | (~a3 | (r | u)),
  \[9]  = (a & (~u & (s & ~r))) | ((a & (~u & (~r & i))) | ((a & (u & (s & r))) | ((a & (u & (r & i))) | ((~u & (~s & (~r & i))) | ((u & (~s & (r & i))) | ((a & (s & ~q)) | ((a & (~q & i)) | ((~u & (~r & q)) | ((u & (r & q)) | (~s & (~q & i))))))))))),
  z1 = (~s & (~q & ~k)) | ((s & (~q & ~c)) | (~q & (~k & ~c))),
  z2 = (~s & (~q & ~p)) | ((s & (~q & ~h)) | (~q & (~p & ~h))),
  a2 = ~v & (~w & \x ),
  a3 = ~v & ~w,
  b3 = ~\x  & (~y & (~z & ~a0)),
  c2 = r | (u | (v | w)),
  c3 = ~u | (v | (w | \x )),
  d0 = \[0] ,
  d2 = (~s & (~q & ~l)) | ((s & (~q & ~d)) | (~q & (~l & ~d))),
  d3 = y | (z | (a0 | b0)),
  e0 = \[1] ,
  e2 = ~v & (~w & (~\x  & y)),
  f0 = \[2] ;
endmodule

