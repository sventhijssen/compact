// IWLS benchmark module "cu" printed on Wed May 29 16:07:22 2002
module cu(a, b, c, d, e, f, g, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, \x , y, z);
input
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  i,
  j,
  k,
  l,
  m,
  n,
  o;
output
  p,
  q,
  r,
  s,
  t,
  u,
  v,
  w,
  \x ,
  y,
  z;
wire
  \[7] ,
  \[8] ,
  \[9] ,
  \[10] ,
  \[0] ,
  \[11] ,
  \[1] ,
  \[12] ,
  \[2] ,
  \[3] ,
  \[4] ,
  a1,
  \[5] ,
  \[6] ;
assign
  \[7]  = \[12]  & f,
  \[8]  = (\[11]  & (~\[1]  & (o & (~n & f)))) | (\[12]  & ~f),
  \[9]  = g & o,
  \[10]  = (g & (~f & ~d)) | (\[11]  & g),
  \[0]  = ~\[1] ,
  \[11]  = ~d & ~c,
  \[1]  = (~f & (e & (~d & c))) | (\[11]  & (f & ~e)),
  \[12]  = \[1]  & ~o,
  p = \[0] ,
  q = \[1] ,
  r = \[2] ,
  s = \[3] ,
  t = \[4] ,
  \[2]  = \[7]  & (~b & ~a),
  u = \[5] ,
  v = \[6] ,
  w = \[7] ,
  \x  = \[8] ,
  y = \[9] ,
  z = \[10] ,
  \[3]  = \[7]  & (~\[5]  & a),
  \[4]  = \[7]  & (~\[5]  & b),
  a1 = (m & (b & a)) | ((l & (b & ~a)) | ((k & (~b & a)) | ((j & (~b & ~a)) | (~o | (n | (i | ~f)))))),
  \[5]  = \[7]  & (b & a),
  \[6]  = (\[11]  & (~a1 & e)) | (\[12]  & ~f);
endmodule

