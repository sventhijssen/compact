// IWLS benchmark module "k2" printed on Wed May 29 16:08:51 2002
module k2(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, \x , y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2, b2, c2, d2, e2, f2, g2, h2, i2, j2, k2, l2);
input
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  t,
  u,
  v,
  w,
  \x ,
  y,
  z,
  a0,
  b0,
  c0,
  d0,
  e0,
  f0,
  g0,
  h0,
  i0,
  j0,
  k0,
  l0,
  m0,
  n0,
  o0,
  p0,
  q0,
  r0,
  s0;
output
  z0,
  z1,
  a1,
  a2,
  b1,
  b2,
  c1,
  c2,
  d1,
  d2,
  e1,
  e2,
  f1,
  f2,
  g1,
  g2,
  h1,
  h2,
  i1,
  i2,
  j1,
  j2,
  k1,
  k2,
  l1,
  l2,
  m1,
  n1,
  o1,
  p1,
  q1,
  r1,
  s1,
  t0,
  t1,
  u0,
  u1,
  v0,
  v1,
  w0,
  w1,
  x0,
  x1,
  y0,
  y1;
wire
  z5,
  z6,
  z7,
  j10,
  z8,
  j11,
  z9,
  j12,
  r10,
  r11,
  r12,
  z10,
  z11,
  \[0] ,
  \[1] ,
  c10,
  c11,
  c12,
  \[2] ,
  \[3] ,
  \[4] ,
  k10,
  k11,
  k12,
  \[5] ,
  \[6] ,
  \[7] ,
  s10,
  s11,
  s12,
  \[8] ,
  \[9] ,
  d10,
  d11,
  d12,
  l10,
  l11,
  l12,
  t10,
  t11,
  t12,
  \[10] ,
  e10,
  e11,
  e12,
  \[11] ,
  \[12] ,
  \[13] ,
  m10,
  m11,
  m12,
  \[14] ,
  \[15] ,
  \[16] ,
  u10,
  u11,
  u12,
  \[17] ,
  \[18] ,
  \[19] ,
  \[20] ,
  f10,
  f11,
  f12,
  \[21] ,
  \[22] ,
  \[23] ,
  n10,
  n11,
  n12,
  \[25] ,
  \[26] ,
  v10,
  v11,
  v12,
  \[27] ,
  \[28] ,
  \[29] ,
  \[30] ,
  g10,
  g11,
  g12,
  \[31] ,
  \[32] ,
  \[33] ,
  o10,
  o11,
  o12,
  \[34] ,
  \[35] ,
  \[36] ,
  w10,
  w11,
  \[37] ,
  \[38] ,
  \[39] ,
  \[40] ,
  h10,
  h11,
  h12,
  \[41] ,
  \[42] ,
  \[43] ,
  p10,
  p11,
  p12,
  x10,
  x11,
  a6,
  a7,
  a8,
  a9,
  b6,
  b7,
  b8,
  b9,
  c6,
  c7,
  c8,
  c9,
  d5,
  d6,
  d7,
  d8,
  d9,
  e6,
  e7,
  e8,
  e9,
  f6,
  f7,
  f8,
  f9,
  a10,
  a11,
  g6,
  a12,
  g7,
  g8,
  g9,
  h6,
  h7,
  h8,
  h9,
  i6,
  i7,
  i8,
  i9,
  j6,
  j7,
  i10,
  j8,
  i11,
  j9,
  i12,
  k6,
  k7,
  k8,
  k9,
  l6,
  l7,
  l8,
  l9,
  m6,
  m7,
  m8,
  m9,
  q10,
  q11,
  q12,
  n6,
  n7,
  n8,
  n9,
  o6,
  o7,
  o8,
  o9,
  p6,
  p7,
  p8,
  p9,
  y10,
  y11,
  q6,
  q7,
  q8,
  q9,
  r6,
  r7,
  r8,
  r9,
  s6,
  s7,
  s8,
  s9,
  t6,
  t7,
  t8,
  t9,
  u6,
  u7,
  u8,
  u9,
  v6,
  v7,
  v8,
  v9,
  b10,
  b11,
  w6,
  b12,
  w7,
  w8,
  w9,
  x5,
  x6,
  x7,
  x8,
  x9,
  y5,
  y6,
  y7,
  y8,
  y9;
assign
  z0 = \[6] ,
  z1 = \[32] ,
  z5 = e0 & (~d0 & (c0 & (a0 & (~v & (~u & (t & (s & (~l & a)))))))),
  z6 = e0 & (z & (~v & (~u & (~t & (s & ~k))))),
  z7 = n0 & (~h0 & (~f0 & (e0 & (~d0 & (~c0 & (w & (v & (~u & (~t & (~s & j)))))))))),
  j10 = e0 & (~d0 & (c0 & (v & (~u & (~t & s))))),
  z8 = z & (v & (u & (~t & (~s & ~k)))),
  j11 = ~e0 & (~d0 & (c0 & (~v & (u & (~t & ~s))))),
  z9 = e0 & (d0 & (~c0 & (w & (v & (u & (t & ~s)))))),
  j12 = e0 & (~d0 & (~c0 & (w & (~v & (u & (t & ~s)))))),
  r10 = e0 & (~d0 & (~c0 & (z & (v & (u & (~t & (s & (~k & f)))))))),
  r11 = e0 & (d0 & (c0 & (w & (~v & (u & (t & ~s)))))),
  r12 = ~e0 & (~d0 & (c0 & (w & (~v & (u & (t & ~s)))))),
  z10 = e0 & (~d0 & (~c0 & (z & (v & (u & (~t & (s & (~p & (l & (k & (~f & a))))))))))),
  z11 = e0 & (~d0 & (y & (~v & (u & (~t & ~s))))),
  \[0]  = l11 | (e10 | (n9 | (m9 | (l6 | g9)))),
  \[1]  = l11 | g9,
  c10 = ~e0 & (d0 & (~c0 & (~v & (~u & (~t & (~s & d)))))),
  c11 = e0 & (~d0 & (~c0 & (a0 & (v & (u & (~t & (s & (~p & (~l & (~f & a)))))))))),
  c12 = e0 & (~d0 & (~c0 & (\x  & (~v & (u & (~t & ~s)))))),
  \[2]  = 0,
  \[3]  = n9 | m9,
  \[4]  = l11 | (n9 | l6),
  k10 = e0 & (~d0 & (~c0 & (w & (v & (u & (~t & (s & (~p & (~f & a))))))))),
  k11 = e0 & (z & (v & (~u & (t & (s & ~k))))),
  k12 = e0 & (~d0 & (c0 & (~v & (u & (~t & (~s & (~d & (~c & a)))))))),
  \[5]  = t10 | (f10 | (m6 | h9)),
  \[6]  = g8 | (j8 | (n8 | (z5 | (a6 | (b6 | (e6 | (p6 | (k6 | (s6 | (q6 | (q12 | (u6 | (s11 | (v12 | (k12 | (d12 | (x11 | (t11 | (f11 | (c11 | (z10 | (w10 | (k10 | (\[41]  | (d9 | (c9 | (b9 | (a9 | w8)))))))))))))))))))))))))))),
  \[7]  = e6 | (p6 | (z10 | (w10 | (b9 | a9)))),
  s10 = e0 & (~d0 & (~c0 & (z & (v & (u & (~t & (s & (~p & (~k & (~f & a)))))))))),
  s11 = ~e0 & (d0 & (c0 & (w & (~v & (u & (t & (~s & a))))))),
  s12 = e0 & (~d0 & (~c0 & (a0 & (~v & (u & (t & ~s)))))),
  \[8]  = j8 | (z5 | (e6 | (k6 | (s6 | (s11 | (k12 | (t11 | (c11 | (w10 | (k10 | (\[41]  | (c9 | (a9 | w8))))))))))))),
  \[9]  = g8 | (d12 | x11),
  d10 = ~e0 & (d0 & (~c0 & (~v & (~u & (~t & (~s & (f & ~d))))))),
  d11 = ~e0 & (d0 & (~c0 & (a0 & (v & (u & (~t & (s & ~l))))))),
  d12 = ~e0 & (d0 & (~c0 & (\x  & (~v & (u & (~t & (~s & a))))))),
  l10 = ~e0 & (d0 & (~c0 & (w & (v & (u & (~t & s)))))),
  l11 = e0 & (~d0 & (y & (v & (u & (t & (s & ~a)))))),
  l12 = ~e0 & (d0 & (c0 & (~v & (u & (~t & ~s))))),
  t10 = e0 & (~d0 & (v & (u & (t & (s & a))))),
  t11 = ~e0 & (d0 & (~c0 & (~v & (~u & (~t & (~s & (~f & (~d & a)))))))),
  t12 = ~e0 & (d0 & (~c0 & (w & (~v & (u & (t & (~s & f))))))),
  \[10]  = q7 | (t7 | (u7 | (v7 | (w7 | (x7 | (y7 | (z7 | (d8 | (f8 | (i8 | (m8 | (y5 | (f6 | (g6 | (j6 | (\[21]  | (\[20]  | (g12 | (r11 | (u12 | (i12 | (n12 | (l12 | (d7 | (y11 | (u11 | (x9 | (h11 | (g11 | (e11 | (d11 | (a11 | (x10 | (l10 | (g10 | (y9 | (o6 | (p9 | (o9 | (i9 | (f9 | (e9 | x8)))))))))))))))))))))))))))))))))))))))))),
  e10 = e0 & (~d0 & (~c0 & (v & (~u & (~t & (s & ~a)))))),
  e11 = e0 & (d0 & (~c0 & (a0 & (v & (u & (~t & (s & ~l))))))),
  e12 = e0 & (~d0 & (~c0 & (~b0 & (~v & (u & (t & s)))))),
  \[11]  = o7 | (f8 | (h8 | (m8 | (d6 | (f6 | (r6 | (g12 | (u12 | (l12 | (d7 | (y11 | (u11 | (x9 | (h11 | (g11 | (e11 | (d11 | (b11 | (y10 | (x10 | (m10 | (l10 | (h10 | (g10 | (z9 | (y9 | (t6 | (o6 | (s9 | (r9 | (p9 | (o9 | (j9 | (i9 | (f9 | (e9 | (y8 | x8))))))))))))))))))))))))))))))))))))),
  \[12]  = p7 | (q7 | (d8 | (f8 | (h8 | (i8 | (m8 | (y5 | (d6 | (f6 | (g6 | (j6 | (\[21]  | (\[20]  | (r6 | (g12 | (r11 | (u12 | (i12 | (n12 | (l12 | (d7 | (y11 | (u11 | (b10 | (x9 | (t9 | (l9 | (h11 | (g11 | (e11 | (d11 | (b11 | (a11 | (y10 | (x10 | (m10 | (l10 | (h10 | (g10 | (z9 | (y9 | (t6 | (o6 | (s9 | (r9 | (j9 | (i9 | (f9 | (e9 | (y8 | x8)))))))))))))))))))))))))))))))))))))))))))))))))),
  \[13]  = q7 | (t7 | (u7 | (v7 | (w7 | (z7 | (h8 | (i8 | (e12 | (y5 | (d6 | (c6 | (g6 | (h6 | (j6 | (n6 | (\[21]  | (\[20]  | (r6 | (v6 | (w6 | (x6 | (y6 | (o11 | (r11 | (o12 | (s12 | (p12 | (j12 | (i12 | (v10 | (n12 | (m12 | (c12 | (p11 | (b10 | (t9 | (l9 | (a11 | (p9 | (o9 | (u8 | r8))))))))))))))))))))))))))))))))))))))))),
  m10 = e0 & (d0 & (~c0 & (w & (v & (u & (~t & s)))))),
  m11 = e0 & (w & (v & (u & (t & s)))),
  m12 = e0 & (~d0 & (w & (~v & (~u & (t & ~s))))),
  \[14]  = r7 | (t7 | (v7 | (x7 | (z7 | (c8 | (h8 | (i8 | (y5 | (d6 | (g6 | (j6 | (\[21]  | (\[20]  | (r6 | (o11 | (r11 | (o12 | (i12 | (n12 | (t9 | (h11 | (e11 | (a11 | (z9 | (t6 | (p9 | f9)))))))))))))))))))))))))),
  \[15]  = g7 | (i7 | (j7 | (l7 | (m7 | (n7 | (o7 | (s7 | (e8 | (f8 | (g8 | (i8 | (k8 | (m8 | (o8 | (y5 | (f6 | (c6 | (g6 | (j6 | (\[21]  | (\[20]  | (g12 | (w6 | (u9 | (r11 | (u12 | (t12 | (i12 | (n12 | (m12 | (l12 | (k12 | (f12 | (q11 | (d7 | (z11 | (y11 | (x11 | (u11 | (d10 | (c10 | (x9 | (g11 | (d11 | (a11 | (x10 | (l10 | (i10 | (g10 | (f10 | (y9 | (o6 | (p9 | (o9 | (i9 | (e9 | (x8 | (u8 | r8)))))))))))))))))))))))))))))))))))))))))))))))))))))))))),
  \[16]  = q7 | (t7 | (u7 | (v7 | (w7 | (x7 | (y7 | (z7 | (d8 | (e8 | (g8 | (h8 | (i8 | (k8 | (m8 | (o8 | (q8 | (e12 | (y5 | (d6 | (c6 | (g6 | (h6 | (j6 | (n6 | (\[21]  | (\[20]  | (r6 | (v6 | (w6 | (y6 | (u9 | (o11 | (r11 | (o12 | (t12 | (s12 | (p12 | (i12 | (n12 | (k12 | (f12 | (q11 | (a12 | (d5 | (x11 | (d10 | (c10 | (g11 | (d11 | (a11 | (e9 | (u8 | r8)))))))))))))))))))))))))))))))))))))))))))))))))))),
  u10 = c0 & (v & (u & (~t & (s & (~q & h))))),
  u11 = e0 & (d0 & (~c0 & (~v & (~u & (~t & ~s))))),
  u12 = e0 & (d0 & (~c0 & (w & (~v & (u & (t & ~s)))))),
  \[17]  = g7 | (h7 | (n7 | (o7 | (p7 | (r7 | (s7 | (c8 | (e8 | (f8 | (i8 | (q8 | (y5 | (d6 | (f6 | (c6 | (g6 | (j6 | (\[21]  | (\[20]  | (r6 | (g12 | (w6 | (x6 | (y6 | (o11 | (r11 | (o12 | (u12 | (p12 | (m12 | (l12 | (d7 | (z11 | (y11 | (u11 | (b10 | (x9 | (t9 | (l9 | (i11 | (h11 | (e11 | (b11 | (a11 | (y10 | (x10 | (m10 | (l10 | (j10 | (h10 | (g10 | (z9 | (y9 | (t6 | (o6 | (s9 | (r9 | (p9 | (o9 | (j9 | (i9 | (f9 | (e9 | (y8 | (x8 | (u8 | r8)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))),
  \[18]  = g7 | (h7 | (i7 | (j7 | (e8 | (f8 | (h8 | (e12 | (f6 | (h6 | (n6 | (g12 | (v6 | (y6 | (b7 | (u12 | (s12 | (p12 | (j12 | (i12 | (v10 | (n12 | (m12 | (l12 | (d7 | (c12 | (z11 | (y11 | (u11 | (p11 | (x9 | (x10 | (l10 | (j10 | (g10 | (f10 | (y9 | (o6 | (p9 | (o9 | (i9 | (x8 | (u8 | r8)))))))))))))))))))))))))))))))))))))))))),
  \[19]  = i7 | (k7 | (l7 | (o7 | (s7 | (e8 | (f8 | (h8 | (m8 | (e12 | (d6 | (f6 | (c6 | (h6 | (n6 | (r6 | (g12 | (v6 | (w6 | (x6 | (o11 | (o12 | (u12 | (p12 | (j12 | (i12 | (v10 | (m12 | (l12 | (d7 | (c12 | (a12 | (d5 | (y11 | (u11 | (p11 | (x9 | (g11 | (d11 | (x10 | (l10 | (g10 | (f10 | (y9 | (o6 | (p9 | (o9 | (i9 | (e9 | x8)))))))))))))))))))))))))))))))))))))))))))))))),
  \[20]  = e0 & (d0 & (~c0 & (a0 & (~v & (u & (~t & (s & ~r))))))),
  f10 = e0 & (~d0 & (~c0 & (v & (~u & (~t & (s & a)))))),
  f11 = e0 & (~d0 & (~c0 & (a0 & (v & (u & (~t & (s & (~p & (l & (~f & a)))))))))),
  f12 = e0 & (~d0 & (c0 & (~v & (u & (~t & (~s & (g & (~d & ~c)))))))),
  \[21]  = ~e0 & (d0 & (c0 & (a0 & (~v & (u & (~t & s)))))),
  \[22]  = g7 | (h7 | (i7 | (j7 | (k7 | (l7 | (m7 | (n7 | (o7 | (p7 | (q7 | (r7 | (s7 | (t7 | (u7 | (v7 | (w7 | (x7 | (y7 | (z7 | (c8 | (d8 | (e8 | (f8 | (g8 | (h8 | (i8 | (k8 | (m8 | (o8 | (q8 | (e12 | (y5 | (d6 | (f6 | (c6 | (g6 | (h6 | (i6 | (j6 | (n6 | (\[21]  | (\[20]  | (r6 | (g12 | (v6 | (w6 | (x6 | (y6 | (z6 | (b7 | (u9 | (o11 | (r11 | (o12 | (u12 | (t12 | (s12 | (p12 | (j12 | (i12 | (v10 | (n12 | (m12 | (k12 | (f12 | (q11 | (d7 | (c12 | (a12 | (z11 | (d5 | (x11 | (u11 | (d10 | (c10 | (p11 | (b10 | (x9 | (k11 | (t9 | (l9 | (i11 | (h11 | (g11 | (e11 | (d11 | (b11 | (a11 | (y10 | (x10 | (s10 | (r10 | (m10 | (l10 | (j10 | (i10 | (h10 | (g10 | (f10 | (z9 | (y9 | (t6 | (o6 | (s9 | (r9 | (q9 | (p9 | (o9 | (j9 | (i9 | (f9 | (e9 | (z8 | (y8 | (x8 | r8))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))),
  \[23]  = g11 | (d11 | e9),
  n10 = e0 & (~d0 & (~c0 & (v & (u & (~t & (s & (p & ~f))))))),
  n11 = e0 & (~d0 & (c0 & (~v & (u & (~t & (~s & (~g & (~d & ~c)))))))),
  n12 = ~e0 & (d0 & (w & (~v & (~u & (t & (~s & b)))))),
  \[25]  = n7 | (e12 | (c6 | (h6 | (i6 | (n6 | (v6 | (w6 | (x6 | (y6 | (z6 | (b7 | (q10 | (s12 | (p12 | (j12 | (v10 | (m12 | (c12 | (b12 | (z11 | (d5 | (p11 | (m11 | (k11 | (s10 | (r10 | (q9 | (z8 | u8)))))))))))))))))))))))))))),
  \[26]  = e12 | (j12 | (c12 | p11)),
  v10 = e0 & (~d0 & (\x  & (~v & (~u & (t & ~s))))),
  v11 = ~e0 & (~d0 & (c0 & (~v & (~u & (~t & ~s))))),
  v12 = ~e0 & (d0 & (~c0 & (w & (~v & (u & (t & (~s & (~f & a)))))))),
  \[27]  = g8 | (k8 | (o8 | (u9 | (t12 | (k12 | (f12 | (q11 | (x11 | (d10 | c10))))))))),
  \[28]  = f7 | (g7 | (h7 | (i7 | (j7 | (k7 | (l7 | (m7 | (p7 | (s7 | (z6 | (b7 | (q10 | (b12 | (a12 | (d5 | (b10 | (m11 | (k11 | (t9 | (l9 | (i11 | (h11 | (b11 | (u10 | (e7 | (s10 | (r10 | (x5 | (p10 | (j10 | (k9 | (a7 | (v9 | (t6 | (s9 | (r9 | (q9 | (j9 | (f9 | (z8 | y8)))))))))))))))))))))))))))))))))))))))),
  \[29]  = g8 | (n8 | (b6 | (u6 | (v12 | (k12 | (d12 | (x11 | (t11 | (t10 | (f11 | (c11 | (z10 | (w10 | (k10 | (f10 | (\[41]  | (m6 | (h9 | (d9 | (c9 | (b9 | (a9 | w8)))))))))))))))))))))),
  \[30]  = j8 | (e6 | (p6 | (k6 | (q12 | s11)))),
  g10 = ~e0 & (d0 & (~c0 & (v & (~u & (~t & s))))),
  g11 = ~e0 & (d0 & (~c0 & (a0 & (v & (u & (~t & (s & l))))))),
  g12 = ~e0 & (d0 & (~c0 & (a0 & (~v & (u & (~t & (s & r))))))),
  \[31]  = j8 | (z5 | (a6 | (s6 | (q6 | s11)))),
  \[32]  = ~e0 & (~d0 & (~c0 & (~b0 & (v & (~o & (~n & ~m)))))),
  \[33]  = f8 | (g8 | (i8 | (k8 | o8))),
  o10 = c0 & (v & (u & (~t & (s & (~q & ~h))))),
  o11 = e0 & (~d0 & (c0 & (w & (~v & (u & (t & (~s & (~d & ~c)))))))),
  o12 = e0 & (~d0 & (c0 & (w & (~v & (u & (t & (~s & d))))))),
  \[34]  = o7 | (q7 | (r7 | (t7 | (v7 | (w7 | (x7 | (y7 | (z7 | (a8 | (b8 | (c8 | (j8 | (l8 | (m8 | (n8 | (z5 | (a6 | (d6 | (f6 | (s6 | (q6 | (r6 | (g12 | (o11 | (s11 | (o12 | (r12 | (u12 | (k12 | (j11 | (d7 | (x11 | (v11 | (u11 | (e11 | (y10 | (m10 | (i10 | (h10 | (z9 | (o6 | (m6 | (n9 | (m9 | l6)))))))))))))))))))))))))))))))))))))))))))),
  \[35]  = n7 | (u7 | (d8 | (f8 | (h8 | (j8 | (k8 | (l8 | (o8 | (q8 | (e12 | (z5 | (a6 | (b6 | (c6 | (e6 | (p6 | (h6 | (k6 | (n6 | (s6 | (q6 | (q12 | (u6 | (v6 | (w6 | (o11 | (r11 | (s11 | (o12 | (v12 | (j12 | (v10 | (m12 | (k12 | (n11 | (h12 | (d12 | (c12 | (z11 | (x11 | (w11 | (t11 | (p11 | (x9 | (t10 | (g11 | (f11 | (d11 | (c11 | (a11 | (z10 | (x10 | (w10 | (l10 | (k10 | (g10 | (f10 | (y9 | (\[41]  | (o6 | (m6 | (p9 | (o9 | (i9 | (h9 | (e9 | (d9 | (c9 | (b9 | (a9 | (x8 | w8))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))),
  \[36]  = r7 | (u7 | (c8 | (g8 | (h8 | (j8 | (m8 | (q8 | (d6 | (b6 | (e6 | (p6 | (k6 | (r6 | (q12 | (u6 | (s11 | (r12 | (v12 | (j11 | (d12 | (v11 | (t11 | (x9 | (g11 | (d11 | (a11 | (y10 | (x10 | (p8 | (o10 | (n10 | (l10 | (i10 | (g10 | (c7 | (a10 | (y9 | (w9 | (o6 | (n9 | (m9 | (l6 | (i9 | (e9 | (x8 | (\[32]  | (v8 | (t8 | s8)))))))))))))))))))))))))))))))))))))))))))))))),
  w10 = e0 & (~d0 & (~c0 & (z & (v & (u & (~t & (s & (~p & (~l & (k & (~f & a))))))))))),
  w11 = e0 & (~d0 & (c0 & (~v & (~u & (~t & (~s & (~d & ~c))))))),
  \[37]  = (e0 & (a0 & (v & (u & (t & s))))) | (f7 | (g7 | (h7 | (i7 | (j7 | (k7 | (l7 | (m7 | (n7 | (o7 | (p7 | (q7 | (r7 | (s7 | (t7 | (u7 | (v7 | (w7 | (x7 | (y7 | (z7 | (a8 | (b8 | (c8 | (d8 | (e8 | (f8 | (g8 | (h8 | (i8 | (j8 | (k8 | (l8 | (m8 | (n8 | (o8 | (q8 | (e12 | (y5 | (z5 | (a6 | (d6 | (f6 | (b6 | (c6 | (g6 | (e6 | (p6 | (h6 | (i6 | (j6 | (k6 | (n6 | (\[21]  | (s6 | (q6 | (\[20]  | (r6 | (q12 | (g12 | (u6 | (v6 | (w6 | (x6 | (y6 | (z6 | (b7 | (q10 | (u9 | (o11 | (r11 | (s11 | (o12 | (r12 | (u12 | (v12 | (t12 | (s12 | (p12 | (j12 | (i12 | (v10 | (n12 | (m12 | (l12 | (k12 | (f12 | (q11 | (n11 | (h12 | (j11 | (d7 | (d12 | (c12 | (b12 | (a12 | (z11 | (d5 | (y11 | (x11 | (w11 | (v11 | (u11 | (t11 | (d10 | (c10 | (p11 | (b10 | (x9 | (t10 | (m11 | (k11 | (t9 | (l9 | (i11 | (h11 | (g11 | (f11 | (e11 | (d11 | (c11 | (b11 | (a11 | (z10 | (y10 | (x10 | (w10 | (p8 | (u10 | (e7 | (s10 | (r10 | (x5 | (p10 | (o10 | (n10 | (m10 | (l10 | (k10 | (j10 | (i10 | (h10 | (g10 | (f10 | (k9 | (c7 | (a7 | (a10 | (z9 | (y9 | (\[41]  | (w9 | (v9 | (t6 | (o6 | (m6 | (s9 | (r9 | (q9 | (p9 | (o9 | (n9 | (m9 | (l6 | (j9 | (i9 | (h9 | (f9 | (e9 | (d9 | (c9 | (b9 | (a9 | (z8 | (y8 | (x8 | (w8 | (\[32]  | (v8 | (t8 | (s8 | r8))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))),
  \[38]  = (~p & (~f & (~a & (e0 & (~d0 & (~c0 & (w & (v & (u & (t & ~s)))))))))) | ((~c & (~d & (~a & (e0 & (~d0 & (c0 & (~v & (~u & (~t & ~s))))))))) | ((c & (~d & (~a & (e0 & (~d0 & (c0 & (~v & (u & (~t & ~s))))))))) | ((~p & (~f & (~a & (e0 & (~d0 & (~c0 & (v & (u & (~t & s))))))))) | ((~f & (~b0 & (~a & (e0 & (d0 & (~c0 & (~v & (u & (t & s))))))))) | ((~f & (~d & (~a & (~e0 & (d0 & (~c0 & (~v & (~u & (~t & ~s))))))))) | ((~f & (~a & (~e0 & (d0 & (~c0 & (w & (~v & (u & (t & ~s))))))))) | ((~e & (~b0 & (~a & (~e0 & (d0 & (c0 & (~v & (u & (t & s))))))))) | ((~r & (a0 & (~a & (~e0 & (d0 & (~c0 & (~v & (u & (~t & s))))))))) | ((r & (a0 & (~a & (~e0 & (d0 & (~c0 & (~v & (u & (~t & s))))))))) | ((l & (a0 & (~a & (e0 & (~d0 & (c0 & (~v & (u & (~t & s))))))))) | ((\x  & (~a & (~e0 & (d0 & (~c0 & (~v & (u & (~t & ~s)))))))) | ((\x  & (e0 & (~d0 & (~c0 & (v & (~u & (t & (~s & ~b)))))))) | ((a0 & (~a & (~e0 & (d0 & (~c0 & (~v & (~u & (t & s)))))))) | ((a0 & (~a & (e0 & (~d0 & (c0 & (~v & (~u & (t & s)))))))) | ((~a & (~e0 & (d0 & (c0 & (w & (~v & (u & (t & ~s)))))))) | ((e0 & (~d0 & (~c0 & (w & (v & (~u & (t & (~s & ~b)))))))) | ((\x  & (~e0 & (d0 & (~v & (~u & (t & (~s & ~b))))))) | ((b0 & (d & (~a & (~d0 & (~v & (u & (t & s))))))) | ((z & (~a & (~e0 & (d0 & (~v & (~u & (t & s))))))) | ((z & (~a & (e0 & (~d0 & (v & (u & (~t & ~s))))))) | ((a0 & (~a & (e0 & (~d0 & (v & (u & (~t & ~s))))))) | ((~a & (~e0 & (d0 & (w & (~v & (~u & (t & s))))))) | ((~a & (e0 & (~d0 & (w & (v & (u & (~t & ~s))))))) | ((~e0 & (d0 & (w & (~v & (~u & (t & (~s & ~b))))))) | ((~a & (e0 & (~d0 & (c0 & (v & (t & ~s)))))) | (l11 | (e10 | g9))))))))))))))))))))))))))),
  \[39]  = f8 | (k8 | (y5 | (g6 | (j6 | (\[21]  | (\[20]  | (u9 | (t12 | (i12 | (n12 | (l12 | (d7 | (y11 | (x9 | (g11 | (d11 | (a11 | (x10 | (l10 | (g10 | (y9 | (o6 | (p9 | (o9 | (i9 | (e9 | x8)))))))))))))))))))))))))),
  \[40]  = o8 | (t12 | (d10 | (c10 | (x5 | (p10 | v9))))),
  h10 = e0 & (d0 & (~c0 & (v & (~u & (~t & s))))),
  h11 = e0 & (d0 & (~c0 & (a0 & (v & (u & (~t & (s & l))))))),
  h12 = e0 & (~d0 & (c0 & (~v & (u & (~t & (~s & (~g & d))))))),
  \[41]  = e0 & (~d0 & (~c0 & (w & (v & (u & (t & (~s & (~p & (~f & a))))))))),
  \[42]  = 0,
  \[43]  = z11 | d5,
  p10 = e0 & (~d0 & (~c0 & (~z & (v & (u & (~t & (s & f))))))),
  p11 = e0 & (~d0 & (~c0 & (~v & (~u & (~t & ~s))))),
  p12 = e0 & (~d0 & (~c0 & (\x  & (~v & (u & (t & ~s)))))),
  x10 = ~e0 & (d0 & (~c0 & (z & (v & (u & (~t & (s & ~l))))))),
  x11 = e0 & (~d0 & (c0 & (~v & (~u & (~t & (~s & (~d & (c & a)))))))),
  a1 = \[7] ,
  a2 = \[33] ,
  a6 = e0 & (~d0 & (c0 & (a0 & (~v & (~u & (t & (s & (l & a)))))))),
  a7 = ~e0 & (~d0 & (c0 & (w & (v & (u & (t & (~s & (q & i)))))))),
  a8 = ~n0 & (~h0 & (~f0 & (e0 & (~d0 & (~c0 & (w & (v & (~u & (~t & (~s & j)))))))))),
  a9 = e0 & (~d0 & (z & (v & (u & (~t & (~s & (~l & (k & a)))))))),
  b1 = \[8] ,
  b2 = \[34] ,
  b6 = ~e0 & (d0 & (~c0 & (a0 & (~v & (~u & (t & (s & a))))))),
  b7 = e0 & (z & (~v & (~u & (~t & (s & k))))),
  b8 = f0 & (e0 & (~d0 & (~c0 & (w & (v & (~u & (~t & (~s & j)))))))),
  b9 = e0 & (~d0 & (z & (v & (u & (~t & (~s & (l & (k & a)))))))),
  c1 = \[9] ,
  c2 = \[35] ,
  c6 = e0 & (~d0 & (~c0 & (a0 & (~v & (~u & (t & s)))))),
  c7 = ~e0 & (~d0 & (c0 & (w & (v & (u & (t & (~s & (~q & ~h)))))))),
  c8 = h0 & (e0 & (~d0 & (~c0 & (w & (v & (~u & (~t & (~s & j)))))))),
  c9 = e0 & (~d0 & (a0 & (v & (u & (~t & (~s & (~l & a))))))),
  d1 = \[10] ,
  d2 = \[36] ,
  d5 = e0 & (~d0 & (w & (~v & (u & (~t & ~s))))),
  d6 = ~e0 & (~d0 & (c0 & (a0 & (~v & (~u & (t & s)))))),
  d7 = e0 & (d0 & (~c0 & (~v & (u & (~t & ~s))))),
  d8 = e0 & (~d0 & (~c0 & (w & (v & (~u & (~t & (~s & ~j))))))),
  d9 = e0 & (~d0 & (a0 & (v & (u & (~t & (~s & (l & a))))))),
  e1 = \[11] ,
  e2 = \[37] ,
  e6 = ~e0 & (d0 & (z & (~v & (~u & (t & (s & (~l & (k & a)))))))),
  e7 = c0 & (v & (u & (~t & (s & (q & i))))),
  e8 = ~e0 & (d0 & (~c0 & (b0 & (~v & (u & (t & s)))))),
  e9 = ~e0 & (d0 & (a0 & (v & (u & (~t & ~s))))),
  f1 = \[12] ,
  f2 = \[38] ,
  f6 = e0 & (d0 & (~c0 & (a0 & (~v & (~u & (t & s)))))),
  f7 = ~l0 & (~k0 & (~j0 & (~i0 & (~h0 & (~g0 & (~f0 & (~e0 & (d0 & (\x  & (v & (~u & (~t & ~s)))))))))))),
  f8 = e0 & (~d0 & (b0 & (~v & (u & (t & s))))),
  f9 = e0 & (d0 & (a0 & (v & (u & (~t & ~s))))),
  g1 = \[13] ,
  g2 = \[39] ,
  a10 = ~e0 & (~d0 & (c0 & (w & (v & (u & (t & (~s & (q & ~i)))))))),
  a11 = ~e0 & (d0 & (~c0 & (z & (v & (u & (~t & (s & l))))))),
  g6 = e0 & (d0 & (z & (~v & (~u & (t & s))))),
  a12 = ~e0 & (d0 & (y & (~v & (u & (~t & ~s))))),
  g7 = l0 & (~k0 & (~j0 & (~i0 & (~h0 & (~g0 & (~f0 & (~e0 & (d0 & (\x  & (v & (~u & (~t & ~s)))))))))))),
  g8 = ~e0 & (~d0 & (b0 & (~v & (u & (t & (s & (d & a))))))),
  g9 = e0 & (~d0 & (y & (v & (u & (~t & (~s & ~a)))))),
  h1 = \[14] ,
  h2 = \[40] ,
  h6 = e0 & (~d0 & (z & (~v & (~u & (t & (s & k)))))),
  h7 = k0 & (~j0 & (~i0 & (~h0 & (~g0 & (~f0 & (~e0 & (d0 & (\x  & (v & (~u & (~t & ~s))))))))))),
  h8 = ~e0 & (~d0 & (b0 & (~v & (u & (t & (s & ~d)))))),
  h9 = e0 & (~d0 & (y & (v & (u & (~t & (~s & a)))))),
  i1 = \[15] ,
  i2 = \[41] ,
  i6 = e0 & (~d0 & (z & (~v & (~u & (t & (s & ~k)))))),
  i7 = j0 & (~i0 & (~h0 & (~g0 & (~f0 & (~e0 & (d0 & (\x  & (v & (~u & (~t & ~s)))))))))),
  i8 = e0 & (d0 & (c0 & (~b0 & (~v & (u & (t & s)))))),
  i9 = ~e0 & (d0 & (y & (v & (u & (~t & ~s))))),
  j1 = \[16] ,
  j2 = \[42] ,
  j6 = e0 & (d0 & (w & (~v & (~u & (t & s))))),
  j7 = i0 & (~h0 & (~g0 & (~f0 & (~e0 & (d0 & (\x  & (v & (~u & (~t & ~s))))))))),
  i10 = ~e0 & (~d0 & (c0 & (v & (~u & (~t & s))))),
  j8 = ~e0 & (d0 & (c0 & (~b0 & (~v & (u & (t & (s & (~e & ~a)))))))),
  i11 = e0 & (w & (v & (~u & (t & s)))),
  j9 = e0 & (d0 & (y & (v & (u & (~t & ~s))))),
  i12 = ~e0 & (d0 & (\x  & (~v & (~u & (t & (~s & b)))))),
  k1 = \[17] ,
  k2 = \[43] ,
  k6 = ~e0 & (d0 & (w & (~v & (~u & (t & (s & a)))))),
  k7 = h0 & (~g0 & (~f0 & (~e0 & (d0 & (\x  & (v & (~u & (~t & ~s)))))))),
  k8 = ~e0 & (d0 & (c0 & (~b0 & (~v & (u & (t & (s & e))))))),
  k9 = ~e0 & (~d0 & (c0 & (w & (v & (u & (t & (~s & (~q & h)))))))),
  l1 = \[18] ,
  l2 = d5,
  l6 = e0 & (~d0 & (~c0 & (y & (v & (t & ~s))))),
  l7 = g0 & (~f0 & (~e0 & (d0 & (\x  & (v & (~u & (~t & ~s))))))),
  l8 = e0 & (~d0 & (c0 & (~b0 & (~v & (u & (t & s)))))),
  l9 = e0 & (z & (v & (~u & (t & (s & k))))),
  m1 = \[19] ,
  m6 = e0 & (~d0 & (c0 & (v & (t & (~s & a))))),
  m7 = f0 & (~e0 & (d0 & (\x  & (v & (~u & (~t & ~s)))))),
  m8 = ~e0 & (~d0 & (c0 & (~b0 & (~v & (u & (t & s)))))),
  m9 = e0 & (~d0 & (~c0 & (z & (v & (t & (~s & k)))))),
  q10 = e0 & (w & (~v & (~u & (~t & s)))),
  q11 = e0 & (~d0 & (c0 & (~v & (u & (~t & (~s & (g & d))))))),
  q12 = ~e0 & (d0 & (~c0 & (a0 & (~v & (u & (~t & (s & (~r & a)))))))),
  n1 = \[20] ,
  n6 = e0 & (~d0 & (w & (~v & (~u & (t & s))))),
  n7 = e0 & (~d0 & (\x  & (v & (~u & (~t & ~s))))),
  n8 = e0 & (d0 & (~c0 & (~b0 & (~v & (u & (t & (s & (~f & a)))))))),
  n9 = e0 & (~d0 & (~c0 & (a0 & (v & (t & ~s))))),
  o1 = \[21] ,
  o6 = ~e0 & (d0 & (c0 & (v & (t & ~s)))),
  o7 = ~s0 & (r0 & (~q0 & (~p0 & (~o0 & (~n0 & (~m0 & (~e0 & (d0 & (~c0 & (w & (v & (~u & (~t & (~s & ~j)))))))))))))),
  o8 = e0 & (d0 & (~c0 & (~b0 & (~v & (u & (t & (s & f))))))),
  o9 = e0 & (~d0 & (~c0 & (w & (v & (~u & (t & (~s & b))))))),
  p1 = \[22] ,
  p6 = ~e0 & (d0 & (z & (~v & (~u & (t & (s & (l & (k & a)))))))),
  p7 = ~s0 & (~r0 & (~q0 & (~p0 & (~o0 & (~n0 & (~m0 & (~e0 & (d0 & (~c0 & (w & (v & (~u & (~t & (~s & ~j)))))))))))))),
  p8 = c0 & (v & (u & (~t & (s & (q & ~i))))),
  p9 = e0 & (~d0 & (~c0 & (\x  & (v & (~u & (t & (~s & b))))))),
  y10 = e0 & (d0 & (~c0 & (z & (v & (u & (~t & (s & ~l))))))),
  y11 = ~e0 & (d0 & (c0 & (~v & (~u & (~t & ~s))))),
  q1 = \[23] ,
  q6 = e0 & (~d0 & (c0 & (a0 & (~v & (u & (~t & (s & (~l & a)))))))),
  q7 = s0 & (~r0 & (~q0 & (~p0 & (~o0 & (~n0 & (~m0 & (~e0 & (d0 & (~c0 & (w & (v & (~u & (~t & (~s & ~j)))))))))))))),
  q8 = ~e0 & (d0 & (~c0 & (~b0 & (~v & (u & (t & s)))))),
  q9 = e0 & (~d0 & (~c0 & (z & (v & (t & (~s & ~k)))))),
  r1 = d5,
  r6 = ~e0 & (~d0 & (c0 & (a0 & (~v & (u & (~t & (s & r))))))),
  r7 = ~q0 & (~p0 & (o0 & (~n0 & (~m0 & (~e0 & (d0 & (~c0 & (w & (v & (~u & (~t & (~s & ~j)))))))))))),
  r8 = ~e0 & (~d0 & (~c0 & (~b0 & o))),
  r9 = ~e0 & (d0 & (~c0 & (w & (v & (~u & (t & ~s)))))),
  s1 = \[25] ,
  s6 = e0 & (~d0 & (c0 & (a0 & (~v & (u & (~t & (s & (l & a)))))))),
  s7 = e0 & (c0 & (w & (v & (~u & (~t & ~s))))),
  s8 = ~e0 & (~d0 & (~c0 & (~b0 & (~\x  & (~v & (u & (~t & (~s & ~o)))))))),
  s9 = ~e0 & (d0 & (~c0 & (\x  & (v & (~u & (t & ~s)))))),
  t0 = \[0] ,
  t1 = \[26] ,
  t6 = e0 & (d0 & (c0 & (v & (t & ~s)))),
  t7 = e0 & (d0 & (~c0 & (w & (v & (~u & (~t & ~s)))))),
  t8 = ~e0 & (~d0 & (~c0 & (~b0 & (~v & (~u & (~t & (s & ~o))))))),
  t9 = e0 & (a0 & (v & (~u & (t & s)))),
  u0 = \[1] ,
  u1 = \[27] ,
  u6 = ~e0 & (d0 & (~c0 & (a0 & (~v & (u & (~t & (s & (r & a)))))))),
  u7 = q0 & (~p0 & (n0 & (~m0 & (~e0 & (d0 & (~c0 & (w & (v & (~u & (~t & (~s & ~j))))))))))),
  u8 = ~e0 & (~d0 & (~c0 & (~b0 & (v & (~o & n))))),
  u9 = e0 & (~d0 & (c0 & (w & (~v & (u & (t & (~s & (~d & c)))))))),
  v0 = \[2] ,
  v1 = \[28] ,
  v6 = e0 & (~d0 & (~c0 & (a0 & (~v & (u & (~t & (s & ~r))))))),
  v7 = ~q0 & (~p0 & (n0 & (~m0 & (~e0 & (d0 & (~c0 & (w & (v & (~u & (~t & (~s & ~j))))))))))),
  v8 = ~e0 & (~d0 & (~c0 & (~b0 & (~v & (~o & n))))),
  v9 = e0 & (~d0 & (~c0 & (w & (v & (u & (t & (~s & f))))))),
  w0 = \[3] ,
  w1 = \[29] ,
  b10 = e0 & (d0 & (v & (u & (t & s)))),
  b11 = e0 & (d0 & (~c0 & (z & (v & (u & (~t & (s & l))))))),
  w6 = e0 & (~d0 & (~c0 & (a0 & (~v & (u & (~t & (s & r))))))),
  b12 = e0 & (~d0 & (a0 & (~v & (u & (~t & ~s))))),
  w7 = q0 & (~p0 & (~n0 & (~m0 & (~e0 & (d0 & (~c0 & (w & (v & (~u & (~t & (~s & ~j))))))))))),
  w8 = e0 & (~d0 & (w & (v & (u & (~t & (~s & a)))))),
  w9 = e0 & (~d0 & (~c0 & (w & (v & (u & (t & (~s & (p & ~f)))))))),
  x0 = \[4] ,
  x1 = \[30] ,
  x5 = e0 & (~d0 & (~c0 & (z & (v & (u & (~t & (s & (k & f)))))))),
  x6 = e0 & (\x  & (~v & (u & (~t & s)))),
  x7 = p0 & (~m0 & (~e0 & (d0 & (~c0 & (w & (v & (~u & (~t & (~s & ~j))))))))),
  x8 = ~e0 & (d0 & (~a0 & (v & (u & (~t & ~s))))),
  x9 = ~e0 & (d0 & (v & (u & (t & s)))),
  y0 = \[5] ,
  y1 = \[31] ,
  y5 = ~e0 & (d0 & (c0 & (a0 & (~v & (~u & (t & s)))))),
  y6 = e0 & (w & (~v & (u & (~t & s)))),
  y7 = m0 & (~e0 & (d0 & (~c0 & (w & (v & (~u & (~t & (~s & ~j)))))))),
  y8 = e0 & (d0 & (~a0 & (v & (u & (~t & ~s))))),
  y9 = ~e0 & (d0 & (~c0 & (w & (v & (u & (t & ~s))))));
endmodule

