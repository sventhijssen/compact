// C7552
module foobar(z6, a7, b7, c7, d7, e7, f7, g7, h7, i7, j7, k7, l7, m7, n7, o7, p7, q7, r7, s7, t7, u7, v7, w7, x7, y7, z7, a8, b8, c8, d8, e8, f8, g8, h8, i8, j8, k8, l8, m8, n8, o8, p8, q8, r8, s8, t8, u8, v8, w8, x8, y8, z8, a9, b9, c9, d9, e9, f9, g9, h9, i9, j9, k9, l9, m9, n9, o9, p9, q9, r9, s9, t9, u9, v9, w9, x9, y9, z9, a10, b10, c10, d10, e10, f10, g10, h10, i10, j10, k10, l10, m10, n10, o10, p10, q10, r10, s10, t10, u10, v10, w10, x10, y10, z10, a11, b11, c11, a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2, b2, c2, d2, e2, f2, g2, h2, i2, j2, k2, l2, m2, n2, o2, p2, q2, r2, s2, t2, u2, v2, w2, x2, y2, z2, a3, b3, c3, d3, e3, f3, g3, h3, i3, j3, k3, l3, m3, n3, o3, p3, q3, r3, s3, t3, u3, v3, w3, x3, y3, z3, a4, b4, c4, d4, e4, f4, g4, h4, i4, j4, k4, l4, m4, n4, o4, p4, q4, r4, s4, t4, u4, v4, w4, x4, y4, z4, a5, b5, c5, d5, e5, f5, g5, h5, i5, j5, k5, l5, m5, n5, o5, p5, q5, r5, s5, t5, u5, v5, w5, x5, y5, z5, a6, b6, c6, d6, e6, f6, g6, h6, i6, j6, k6, l6, m6, n6, o6, p6, q6, r6, s6, t6, u6, v6, w6, x6, y6);
input a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2, b2, c2, d2, e2, f2, g2, h2, i2, j2, k2, l2, m2, n2, o2, p2, q2, r2, s2, t2, u2, v2, w2, x2, y2, z2, a3, b3, c3, d3, e3, f3, g3, h3, i3, j3, k3, l3, m3, n3, o3, p3, q3, r3, s3, t3, u3, v3, w3, x3, y3, z3, a4, b4, c4, d4, e4, f4, g4, h4, i4, j4, k4, l4, m4, n4, o4, p4, q4, r4, s4, t4, u4, v4, w4, x4, y4, z4, a5, b5, c5, d5, e5, f5, g5, h5, i5, j5, k5, l5, m5, n5, o5, p5, q5, r5, s5, t5, u5, v5, w5, x5, y5, z5, a6, b6, c6, d6, e6, f6, g6, h6, i6, j6, k6, l6, m6, n6, o6, p6, q6, r6, s6, t6, u6, v6, w6, x6, y6;
output z6, a7, b7, c7, d7, e7, f7, g7, h7, i7, j7, k7, l7, m7, n7, o7, p7, q7, r7, s7, t7, u7, v7, w7, x7, y7, z7, a8, b8, c8, d8, e8, f8, g8, h8, i8, j8, k8, l8, m8, n8, o8, p8, q8, r8, s8, t8, u8, v8, w8, x8, y8, z8, a9, b9, c9, d9, e9, f9, g9, h9, i9, j9, k9, l9, m9, n9, o9, p9, q9, r9, s9, t9, u9, v9, w9, x9, y9, z9, a10, b10, c10, d10, e10, f10, g10, h10, i10, j10, k10, l10, m10, n10, o10, p10, q10, r10, s10, t10, u10, v10, w10, x10, y10, z10, a11, b11, c11;
not(k8, e);
not(t_0, z15);
not(t_1, n15);
or(o8, t_0, t_1);
not(p8, j15);
not(q8, i15);
not(r8, g15);
not(s8, h15);
not(t_2, x15);
not(t_3, j5);
or(v8, t_2, t_3);
not(w8, u15);
not(t_4, x15);
not(t_5, j5);
or(x8, t_4, t_5);
not(t_6, y15);
not(t_7, k15);
or(y8, t_6, t_7);
not(z8, u15);
not(a9, u18);
and(c9, i2, b9);
not(t_8, o114);
not(t_9, i109);
or(d9, t_8, t_9);
or(e9, v114, a120, z119, b117, n112);
or(f9, k113, l118, k118, m114, y113);
or(g9, i113, n118, m118, n114, y113);
or(h9, u114, v119, u119, c117, l112);
not(t_10, d116);
not(t_11, n119);
or(i9, t_10, t_11);
not(t_12, g116);
not(t_13, o119);
or(j9, t_12, t_13);
not(t_14, j116);
not(t_15, p119);
or(k9, t_14, t_15);
not(t_16, n116);
not(t_17, q119);
or(l9, t_16, t_17);
or(m9, f122, f124);
or(n9, g122, g124);
or(o9, h122, b122);
or(p9, j119, e122);
not(q9, e130);
not(r9, m128);
not(s9, d130);
or(t9, b130, f130);
not(t_18, w126);
not(t_19, g129);
or(u9, t_18, t_19);
not(t_20, l127);
not(t_21, x129);
or(v9, t_20, t_21);
or(w9, f132, o133);
or(x9, h129, u131);
not(t_22, w128);
not(t_23, o131);
or(y9, t_22, t_23);
not(t_24, a129);
not(t_25, r131);
or(z9, t_24, t_25);
not(t_26, c129);
not(t_27, s131);
or(a10, t_26, t_27);
not(t_28, e129);
not(t_29, t131);
or(b10, t_28, t_29);
not(t_30, p129);
not(t_31, z131);
or(c10, t_30, t_31);
not(t_32, t129);
not(t_33, c132);
or(d10, t_32, t_33);
not(t_34, z129);
not(t_35, e132);
or(e10, t_34, t_35);
not(t_36, v129);
not(t_37, d132);
or(f10, t_36, t_37);
not(g10, n133);
or(h10, i129, v131);
or(i10, n128, i131);
or(j10, o128, j131);
or(k10, s128, k131);
or(l10, r128, l131);
not(t_38, f128);
not(t_39, z130);
or(m10, t_38, t_39);
not(t_40, p130);
not(t_41, o132);
or(r10, t_40, t_41);
not(t_42, t130);
not(t_43, r132);
or(s10, t_42, t_43);
not(t_44, v130);
not(t_45, s132);
or(t10, t_44, t_45);
not(t_46, x130);
not(t_47, t132);
or(u10, t_46, t_47);
or(v10, g130, i132);
or(w10, j130, j132);
or(x10, n130, k132);
or(y10, m130, n132);
not(z10, h144);
not(a11, i144);
not(b11, k144);
not(c11, j144);
buf(m13, x6);
buf(n13, x6);
not(o13, w6);
not(p13, v6);
not(q13, u6);
not(r13, t6);
not(s13, s6);
not(t13, r6);
not(u13, q6);
not(v13, p6);
not(w13, o6);
not(x13, n6);
not(y13, m6);
not(z13, l6);
not(a14, k6);
not(b14, j6);
not(c14, i6);
not(d14, h6);
not(e14, g6);
not(f14, f6);
not(g14, e6);
not(h14, d6);
not(i14, c6);
not(j14, c6);
not(k14, b6);
not(l14, b6);
not(m14, a6);
not(n14, z5);
not(o14, y5);
not(p14, y5);
not(q14, x5);
not(r14, w5);
not(s14, v5);
not(t14, u5);
not(u14, t5);
not(v14, s5);
not(w14, r5);
not(t_48, r5);
not(t_49, y6);
or(x14, t_48, t_49);
not(y14, q5);
and(z14, y6, q5);
not(a15, p5);
not(b15, o5);
not(c15, n5);
not(d15, m5);
not(e15, l5);
not(f15, k5);
and(g15, c3, b3, e3, f3);
and(h15, h2, r2, h3, s3);
and(i15, d4, x1, l4, x4);
and(j15, v1, d3, v4, h5);
and(k15, p1, o1);
buf(u8, b1);
not(m15, b1);
not(n15, u);
buf(o15, l);
buf(p15, l);
buf(q15, f);
buf(r15, f);
not(s15, f);
buf(t15, f);
buf(u15, e);
not(t_50, c);
not(t_51, d);
or(v15, t_50, t_51);
not(t_52, c);
not(t_53, d);
or(w15, t_52, t_53);
not(x15, b);
not(y15, b);
not(z15, b);
buf(t8, a);
not(t_54, v14);
not(t_55, y6);
or(b16, t_54, t_55);
and(c16, y6, f15);
not(d16, m13);
not(e16, n13);
buf(f16, o13);
buf(g16, o13);
buf(h16, p13);
buf(i16, p13);
buf(j16, q13);
buf(k16, q13);
buf(l16, r13);
buf(m16, r13);
buf(n16, s13);
buf(o16, s13);
buf(p16, t13);
buf(q16, t13);
buf(r16, u13);
buf(s16, u13);
buf(t16, v13);
buf(u16, v13);
buf(v16, w13);
buf(w16, w13);
buf(x16, y13);
buf(y16, y13);
buf(z16, z13);
buf(a17, z13);
buf(b17, a14);
buf(c17, a14);
buf(d17, b14);
buf(e17, b14);
buf(f17, c14);
buf(g17, c14);
buf(h17, d14);
buf(i17, d14);
buf(j17, e14);
buf(k17, e14);
buf(l17, f14);
buf(m17, f14);
buf(n17, j14);
buf(o17, j14);
buf(p17, l14);
buf(q17, l14);
buf(r17, m14);
buf(s17, m14);
buf(t17, n14);
buf(u17, n14);
buf(v17, p14);
buf(w17, p14);
buf(x17, q14);
buf(y17, q14);
buf(z17, r14);
buf(a18, r14);
buf(b18, s14);
buf(c18, s14);
buf(d18, t14);
buf(e18, t14);
and(f18, x14, p15);
and(g18, x14, p15);
buf(h18, x14);
buf(i18, x14);
not(j18, z14);
buf(k18, a15);
buf(l18, a15);
buf(m18, b15);
buf(n18, b15);
buf(o18, c15);
buf(p18, c15);
buf(q18, d15);
buf(r18, d15);
and(s18, g15, h15);
and(t18, j15, i15);
and(u18, k15, y15);
not(v18, u8);
buf(w18, o15);
buf(x18, o15);
buf(y18, p15);
buf(z18, p15);
buf(a19, p15);
buf(b19, p15);
buf(c19, q15);
buf(d19, q15);
buf(e19, q15);
buf(f19, q15);
not(g19, q15);
buf(h19, r15);
buf(i19, r15);
buf(j19, r15);
buf(k19, r15);
not(l19, r15);
buf(m19, s15);
buf(n19, s15);
buf(o19, t15);
buf(p19, t15);
buf(q19, t15);
buf(r19, t15);
not(s19, t15);
buf(t19, v15);
buf(u19, v15);
buf(v19, v15);
buf(w19, w15);
buf(x19, w15);
buf(y19, w15);
buf(b9, t8);
buf(a20, b16);
not(b20, c16);
not(c20, f16);
not(d20, g16);
not(e20, h16);
not(f20, i16);
not(g20, j16);
not(h20, k16);
not(i20, l16);
not(j20, m16);
not(k20, n16);
not(l20, o16);
not(m20, p16);
not(n20, q16);
not(o20, r16);
not(p20, s16);
not(q20, t16);
not(r20, u16);
not(s20, v16);
not(t20, w16);
not(u20, x16);
not(v20, y16);
not(w20, z16);
not(x20, a17);
not(y20, b17);
not(z20, c17);
not(a21, d17);
not(b21, e17);
not(c21, f17);
not(d21, g17);
not(e21, h17);
not(f21, i17);
not(g21, j17);
not(h21, k17);
not(i21, l17);
not(j21, m17);
and(k21, i14, k19);
not(l21, n17);
not(m21, o17);
and(n21, k14, k19);
not(o21, p17);
not(p21, q17);
and(q21, m14, k19);
not(r21, r17);
not(s21, s17);
not(t21, t17);
not(u21, u17);
and(v21, n14, k19);
and(w21, o14, k19);
not(x21, v17);
not(y21, w17);
not(z21, x17);
not(a22, y17);
and(b22, q14, j19);
and(c22, r14, j19);
not(d22, z17);
not(e22, a18);
not(f22, b18);
not(g22, c18);
and(h22, s14, j19);
not(i22, d18);
and(j22, t14, j19);
not(k22, e18);
and(l22, u14, j19);
and(m22, w14, i19);
not(n22, h18);
not(o22, i18);
and(p22, y14, i19);
buf(q22, j18);
buf(r22, j18);
and(s22, a15, i19);
not(t22, k18);
not(u22, l18);
not(v22, m18);
not(w22, n18);
and(x22, b15, h19);
not(y22, o18);
and(z22, c15, h19);
not(a23, p18);
not(b23, q18);
and(c23, d15, h19);
not(d23, r18);
and(e23, e15, h19);
and(f23, j4, q19);
and(g23, i4, q19);
and(h23, h4, q19);
and(i23, g4, r19);
and(j23, f4, r19);
and(k23, e4, r19);
and(l23, c4, q19);
and(m23, a3, f19);
and(n23, z2, f19);
and(o23, y2, f19);
and(p23, x2, f19);
and(q23, w2, e19);
and(r23, v2, e19);
and(s23, u2, e19);
and(t23, t2, e19);
and(u23, s2, e19);
and(v23, q2, f19);
and(w23, p2, c19);
and(x23, o2, c19);
and(y23, n2, c19);
and(z23, m2, c19);
and(a24, l2, d19);
and(b24, k2, d19);
and(c24, j2, d19);
and(d24, g2, p19);
and(e24, f2, p19);
and(f24, e2, p19);
and(g24, d2, p19);
and(h24, c2, o19);
and(i24, b2, o19);
and(j24, a2, o19);
and(k24, z1, o19);
and(l24, y1, o19);
and(m24, w1, p19);
buf(n24, v18);
buf(o24, v18);
and(p24, m15, h19);
and(q24, d0, m19);
and(r24, p, m19);
and(s24, o, m19);
and(t24, n, n19);
and(u24, m, n19);
not(v24, w18);
and(w24, b16, o15);
not(x24, x18);
and(y24, j18, p15);
and(z24, p15, j18);
not(t_56, p15);
not(t_57, j18);
and(a25, t_56, t_57);
not(b25, y18);
not(c25, z18);
not(t_58, j18);
not(t_59, p15);
and(d25, t_58, t_59);
not(e25, a19);
not(f25, b19);
and(g25, k, m19);
and(h25, j, m19);
and(i25, i, n19);
and(j25, h, n19);
and(k25, g, n19);
not(l25, c19);
not(m25, d19);
not(n25, e19);
not(o25, f19);
buf(p25, g19);
buf(q25, g19);
not(r25, h19);
not(s25, i19);
not(t25, j19);
not(u25, k19);
buf(v25, l19);
buf(w25, l19);
buf(x25, l19);
buf(y25, l19);
not(z25, m19);
not(a26, n19);
not(b26, o19);
not(c26, p19);
not(d26, q19);
not(e26, r19);
buf(f26, s19);
buf(g26, s19);
buf(h26, s19);
buf(i26, s19);
not(t_60, x24);
not(t_61, a20);
or(j26, t_60, t_61);
not(k26, a20);
buf(l26, b20);
and(m26, g14, s25);
and(n26, s5, s25);
not(t_62, c25);
not(t_63, h18);
or(o26, t_62, t_63);
not(t_64, f25);
not(t_65, i18);
or(p26, t_64, t_65);
not(t_66, e25);
not(t_67, q22);
or(q26, t_66, t_67);
not(r26, q22);
not(t_68, b25);
not(t_69, r22);
or(s26, t_68, t_69);
not(t26, r22);
and(u26, k5, s25);
or(v26, f23, d26);
or(w26, g23, d26);
or(x26, h23, d26);
or(y26, i23, e26);
or(z26, j23, e26);
or(a27, k23, e26);
or(b27, l23, d26);
and(c27, b4, a26);
and(d27, a4, a26);
and(e27, z3, a26);
and(f27, y3, a26);
and(g27, r3, a26);
and(h27, m3, z25);
and(i27, l3, z25);
and(j27, k3, z25);
and(k27, j3, z25);
and(l27, i3, z25);
or(m27, q23, n25);
or(n27, r23, n25);
or(o27, s23, n25);
or(p27, t23, n25);
or(q27, u23, n25);
or(r27, w23, l25);
or(s27, x23, l25);
or(t27, y23, l25);
or(u27, z23, l25);
or(v27, a24, m25);
or(w27, b24, m25);
or(x27, c24, m25);
or(y27, h24, b26);
or(z27, i24, b26);
or(a28, j24, b26);
or(b28, k24, b26);
or(c28, l24, b26);
and(d28, u1, c26);
and(e28, u1, o25);
and(f28, t1, c26);
and(g28, t1, o25);
and(h28, s1, o25);
and(i28, s1, c26);
and(j28, r1, c26);
and(k28, r1, o25);
and(l28, q1, c26);
and(m28, q1, o25);
and(n28, n1, p25);
and(o28, n1, f26);
and(p28, m1, f26);
and(q28, m1, p25);
and(r28, l1, f26);
and(s28, l1, p25);
and(t28, k1, g26);
and(u28, k1, q25);
and(v28, j1, q25);
and(w28, j1, g26);
and(x28, i1, q25);
and(y28, i1, g26);
and(z28, h1, r25);
and(a29, g1, r25);
and(b29, f1, r25);
and(c29, e1, r25);
and(d29, d1, u25);
and(e29, c1, u25);
not(f29, n24);
not(g29, o24);
and(h29, a1, p25);
and(i29, a1, f26);
and(j29, z0, f26);
and(k29, z0, p25);
and(l29, y0, g26);
and(m29, y0, q25);
and(n29, x0, g26);
and(o29, x0, q25);
and(p29, v0, s25);
and(q29, u0, r25);
and(r29, t0, u25);
and(s29, s0, t25);
and(t29, r0, t25);
and(u29, q0, t25);
and(v29, p0, t25);
and(w29, o0, x25);
and(x29, n0, y25);
and(y29, m0, y25);
and(z29, l0, x25);
and(a30, k0, x25);
and(b30, j0, v25);
and(c30, i0, v25);
and(d30, h0, v25);
and(e30, g0, w25);
and(f30, f0, v25);
and(g30, f0, s25);
and(h30, e0, v25);
and(i30, d0, i26);
and(j30, c0, t25);
and(k30, b0, u25);
and(l30, a0, u25);
and(m30, z, y25);
and(n30, y, y25);
and(o30, x, y25);
and(p30, w, x25);
and(q30, v, x25);
and(r30, t, w25);
and(s30, s, w25);
and(t30, r, w25);
and(u30, q, w25);
and(v30, p, i26);
and(w30, o, i26);
and(x30, n, h26);
and(y30, m, h26);
and(z30, b20, o15);
buf(a31, y24);
buf(b31, z24);
not(c31, a25);
not(t_70, n22);
not(t_71, z18);
or(d31, t_70, t_71);
not(e31, d25);
not(t_72, o22);
not(t_73, b19);
or(f31, t_72, t_73);
and(g31, k, i26);
and(h31, j, i26);
and(i31, i, h26);
and(j31, h, h26);
and(k31, g, h26);
or(l31, c19, l25);
not(m31, p25);
not(n31, q25);
not(o31, v25);
not(p31, w25);
not(q31, x25);
not(r31, y25);
or(s31, q19, d26);
not(t31, f26);
not(u31, g26);
not(v31, h26);
not(w31, i26);
not(x31, l26);
and(y31, o13, r31);
and(z31, p13, r31);
and(a32, q13, r31);
and(b32, r13, r31);
and(c32, s13, r31);
and(d32, t13, q31);
and(e32, u13, q31);
and(f32, v13, q31);
and(g32, w13, q31);
and(h32, x13, q31);
and(i32, y13, p31);
and(j32, z13, p31);
and(k32, a14, p31);
and(l32, b14, p31);
and(m32, c14, p31);
and(n32, d14, o31);
and(o32, e14, o31);
and(p32, f14, o31);
and(q32, g14, o31);
and(r32, h14, o31);
or(s32, k21, d29);
or(t32, n21, e29);
or(u32, q21, r29);
or(v32, v21, l30);
or(w32, w21, k30);
or(x32, b22, s29);
or(y32, c22, t29);
or(z32, h22, u29);
or(a33, j22, j30);
or(b33, l22, v29);
or(c33, m22, n26);
not(t_74, o26);
not(t_75, d31);
or(d33, t_74, t_75);
not(t_76, p26);
not(t_77, f31);
or(e33, t_76, t_77);
or(f33, p22, u26);
or(g33, s22, p29);
or(h33, x22, b29);
or(i33, z22, c29);
or(j33, c23, a29);
or(k33, e23, z28);
and(l33, g5, v31);
and(m33, f5, v31);
and(n33, e5, v31);
and(o33, d5, v31);
and(p33, c5, t31);
and(q33, b5, t31);
and(r33, a5, t31);
and(s33, z4, t31);
and(t33, y4, t31);
and(u33, w4, v31);
and(v33, u4, u31);
and(w33, t4, u31);
and(x33, s4, u31);
and(y33, r4, u31);
and(z33, q4, w31);
and(a34, p4, w31);
and(b34, o4, w31);
and(c34, n4, w31);
and(d34, m4, w31);
and(e34, k4, u31);
and(f34, x3, m31);
and(g34, w3, m31);
and(h34, v3, m31);
and(i34, u3, m31);
and(j34, t3, m31);
and(k34, q3, n31);
and(l34, p3, n31);
and(m34, o3, n31);
and(n34, n3, n31);
and(o34, g3, n31);
or(p34, m23, h28);
or(q34, n23, k28);
or(r34, o23, g28);
or(s34, p23, m28);
or(t34, v23, e28);
or(u34, d24, i28);
or(v34, e24, j28);
or(w34, f24, f28);
or(x34, g24, l28);
or(y34, m24, d28);
or(z34, p24, q29);
or(a35, q24, l27);
or(b35, r24, k27);
or(c35, s24, h27);
or(d35, t24, c27);
or(e35, u24, g27);
not(t_78, v24);
not(t_79, l26);
or(f35, t_78, t_79);
not(t_80, k26);
not(t_81, x18);
or(g35, t_80, t_81);
not(h35, a31);
not(i35, b31);
not(t_82, t26);
not(t_83, y18);
or(j35, t_82, t_83);
not(t_84, r26);
not(t_85, a19);
or(k35, t_84, t_85);
or(l35, g25, i27);
or(m35, h25, j27);
or(n35, i25, d27);
or(o35, j25, e27);
or(p35, k25, f27);
or(q35, i19, g30);
or(r35, i19, m26);
and(s35, r27, t19);
and(t35, u27, t19);
and(u35, t27, t19);
and(v35, s27, t19);
and(w35, l31, t19);
and(x35, x27, u19);
and(y35, w27, u19);
and(z35, v27, u19);
and(a36, q27, v19);
and(b36, p27, v19);
and(c36, o27, v19);
and(d36, n27, v19);
and(e36, m27, v19);
and(f36, a28, w19);
and(g36, z27, w19);
and(h36, y27, w19);
and(i36, c28, w19);
and(j36, b28, w19);
and(k36, x26, x19);
and(l36, w26, x19);
and(m36, v26, x19);
and(n36, b27, x19);
and(o36, s31, x19);
and(p36, a27, y19);
and(q36, z26, y19);
and(r36, y26, y19);
not(t_86, j26);
not(t_87, g35);
or(s36, t_86, t_87);
and(t36, s32, a36);
buf(u36, s32);
buf(v36, s32);
and(w36, j14, i36);
and(x36, j14, i36);
and(y36, t32, b36);
buf(z36, t32);
buf(a37, t32);
and(b37, l14, j36);
and(c37, l14, j36);
and(d37, m14, f36);
and(e37, m14, f36);
and(f37, u32, c36);
buf(g37, u32);
buf(h37, u32);
and(i37, n14, g36);
and(j37, g36, n14);
not(t_88, g36);
not(t_89, n14);
and(k37, t_88, t_89);
not(t_90, n14);
not(t_91, g36);
and(l37, t_90, t_91);
and(m37, v32, d36);
buf(n37, v32);
buf(o37, v32);
and(p37, w32, e36);
buf(q37, w32);
buf(r37, w32);
and(s37, p14, h36);
and(t37, p14, h36);
and(u37, q14, x34);
and(v37, q14, x34);
and(w37, x32, s34);
buf(x37, x32);
buf(y37, x32);
and(z37, r14, w34);
and(a38, r14, w34);
and(b38, y32, r34);
buf(c38, y32);
buf(d38, y32);
and(e38, s14, v34);
and(f38, s14, v34);
and(g38, z32, q34);
buf(h38, z32);
buf(i38, z32);
and(j38, t14, y34);
and(k38, t14, y34);
not(t_92, t14);
not(t_93, y34);
and(l38, t_92, t_93);
and(m38, a33, t34);
buf(n38, a33);
buf(o38, a33);
not(p38, b33);
not(q38, c33);
buf(r38, d33);
buf(s38, d33);
buf(t38, e33);
buf(u38, e33);
not(v38, f33);
not(t_94, q26);
not(t_95, k35);
or(w38, t_94, t_95);
not(t_96, s26);
not(t_97, j35);
or(x38, t_96, t_97);
and(y38, a15, r36);
and(z38, a15, r36);
and(a39, g33, z35);
buf(b39, g33);
buf(c39, g33);
and(d39, b15, k36);
and(e39, b15, k36);
and(f39, h33, t35);
buf(g39, h33);
buf(h39, h33);
and(i39, c15, m36);
and(j39, c15, m36);
and(k39, i33, v35);
buf(l39, i33);
buf(m39, i33);
and(n39, d15, n36);
and(o39, d15, n36);
not(t_98, d15);
not(t_99, n36);
and(p39, t_98, t_99);
and(q39, j33, w35);
buf(r39, j33);
buf(s39, j33);
not(t39, k33);
not(u39, p34);
buf(v39, q34);
buf(w39, q34);
buf(x39, r34);
buf(y39, r34);
buf(z39, s34);
buf(a40, s34);
buf(b40, t34);
buf(c40, t34);
not(d40, u34);
buf(e40, v34);
buf(f40, v34);
buf(g40, v34);
buf(h40, w34);
buf(i40, w34);
buf(j40, w34);
buf(k40, x34);
buf(l40, x34);
buf(m40, x34);
buf(n40, y34);
buf(o40, y34);
buf(p40, y34);
or(q40, n28, g34);
or(r40, o28, q33);
or(s40, p28, r33);
or(t40, q28, h34);
or(u40, r28, s33);
or(v40, s28, i34);
or(w40, t28, y33);
or(x40, u28, n34);
or(y40, v28, o34);
or(z40, w28, e34);
or(a41, x28, k34);
or(b41, y28, v33);
and(c41, v18, l36);
and(d41, v18, l36);
and(e41, z34, u35);
buf(f41, z34);
buf(g41, z34);
or(h41, h29, f34);
or(i41, i29, p33);
or(j41, j29, t33);
or(k41, k29, j34);
or(l41, l29, w33);
or(m41, m29, l34);
or(n41, n29, x33);
or(o41, o29, m34);
or(p41, w29, d32);
or(q41, x29, c32);
or(r41, y29, b32);
or(s41, z29, f32);
or(t41, a30, g32);
or(u41, b30, o32);
or(v41, c30, n32);
or(w41, d30, p32);
or(x41, e30, m32);
or(y41, f30, q32);
or(z41, h30, r32);
or(a42, i30, d34);
buf(b42, a35);
buf(c42, a35);
or(d42, m30, y31);
or(e42, n30, z31);
or(f42, o30, a32);
or(g42, p30, e32);
or(h42, q30, h32);
or(i42, r30, i32);
or(j42, s30, j32);
or(k42, t30, k32);
or(l42, u30, l32);
or(m42, v30, c34);
buf(n42, b35);
buf(o42, b35);
buf(p42, c35);
buf(q42, c35);
or(r42, w30, z33);
not(s42, d35);
or(t42, x30, l33);
buf(u42, e35);
or(v42, y30, u33);
not(t_100, x31);
not(t_101, w18);
or(w42, t_100, t_101);
and(x42, e33, y24);
and(y42, e33, y24);
and(z42, e33, y24);
and(a43, e33, y24);
and(b43, d33, z24);
buf(c43, l35);
buf(d43, l35);
or(e43, g31, a34);
or(f43, h31, b34);
buf(g43, m35);
buf(h43, m35);
or(i43, i31, m33);
buf(j43, n35);
buf(k43, n35);
or(l43, j31, n33);
buf(m43, o35);
buf(n43, o35);
or(o43, k31, o33);
buf(p43, p35);
buf(q43, p35);
buf(r43, q35);
buf(s43, r35);
buf(t43, r35);
and(u43, s15, e35);
not(v43, s35);
buf(w43, t35);
buf(x43, t35);
buf(y43, u35);
buf(z43, u35);
buf(a44, v35);
buf(b44, v35);
buf(c44, w35);
buf(d44, w35);
not(e44, x35);
not(f44, y35);
buf(g44, z35);
buf(h44, z35);
buf(i44, a36);
buf(j44, a36);
buf(k44, b36);
buf(l44, b36);
buf(m44, c36);
buf(n44, c36);
buf(o44, d36);
buf(p44, d36);
buf(q44, e36);
buf(r44, e36);
buf(s44, f36);
buf(t44, f36);
buf(u44, f36);
buf(v44, g36);
buf(w44, g36);
buf(x44, g36);
buf(y44, h36);
buf(z44, h36);
buf(a45, h36);
buf(b45, i36);
buf(c45, i36);
buf(d45, i36);
buf(e45, j36);
buf(f45, j36);
buf(g45, j36);
buf(h45, k36);
buf(i45, k36);
buf(j45, k36);
buf(k45, l36);
buf(l45, l36);
buf(m45, l36);
buf(n45, m36);
buf(o45, m36);
buf(p45, m36);
buf(q45, n36);
buf(r45, n36);
buf(s45, n36);
not(t45, o36);
not(u45, p36);
not(v45, q36);
buf(w45, r36);
buf(x45, r36);
buf(y45, r36);
and(z45, o13, a42);
and(a46, o13, a42);
and(b46, p13, m42);
and(c46, p13, m42);
and(d46, q13, f43);
and(e46, q13, f43);
and(f46, e43, r13);
and(g46, r13, e43);
not(t_102, r13);
not(t_103, e43);
and(h46, t_102, t_103);
not(t_104, e43);
not(t_105, r13);
and(i46, t_104, t_105);
and(j46, s13, r42);
and(k46, s13, r42);
and(l46, t13, w40);
and(m46, t13, w40);
and(n46, u13, n41);
and(o46, u13, n41);
and(p46, v13, l41);
and(q46, v13, l41);
and(r46, w13, z40);
and(s46, w13, z40);
not(t_106, w13);
not(t_107, z40);
and(t46, t_106, t_107);
and(u46, y13, j41);
and(v46, y13, j41);
and(w46, z13, u40);
and(x46, z13, u40);
and(y46, a14, s40);
and(z46, a14, s40);
and(a47, r40, b14);
and(b47, b14, r40);
not(t_108, b14);
not(t_109, r40);
and(c47, t_108, t_109);
not(t_110, r40);
not(t_111, b14);
and(d47, t_110, t_111);
and(e47, c14, i41);
and(f47, c14, i41);
and(g47, d14, o43);
and(h47, d14, o43);
and(i47, e14, l43);
and(j47, e14, l43);
and(k47, f14, i43);
and(l47, f14, i43);
not(m47, u36);
not(n47, v36);
not(t_112, l21);
not(t_113, c45);
or(o47, t_112, t_113);
not(t_114, m21);
not(t_115, d45);
or(p47, t_114, t_115);
not(q47, z36);
not(r47, a37);
not(t_116, o21);
not(t_117, e45);
or(s47, t_116, t_117);
not(t_118, p21);
not(t_119, f45);
or(t47, t_118, t_119);
not(u47, g37);
not(v47, h37);
not(t_120, r21);
not(t_121, u44);
or(w47, t_120, t_121);
not(t_122, s21);
not(t_123, t44);
or(x47, t_122, t_123);
buf(y47, i37);
buf(z47, j37);
not(t_124, t21);
not(t_125, w44);
or(a48, t_124, t_125);
not(b48, k37);
not(c48, l37);
not(t_126, u21);
not(t_127, v44);
or(d48, t_126, t_127);
not(e48, n37);
not(f48, o37);
not(g48, q37);
not(h48, r37);
not(t_128, x21);
not(t_129, a45);
or(i48, t_128, t_129);
not(t_130, y21);
not(t_131, z44);
or(j48, t_130, t_131);
not(t_132, z21);
not(t_133, m40);
or(k48, t_132, t_133);
not(t_134, a22);
not(t_135, l40);
or(l48, t_134, t_135);
not(m48, x37);
not(n48, y37);
not(o48, c38);
not(p48, d38);
not(t_136, d22);
not(t_137, j40);
or(q48, t_136, t_137);
not(t_138, e22);
not(t_139, i40);
or(r48, t_138, t_139);
not(t_140, f22);
not(t_141, g40);
or(s48, t_140, t_141);
not(t_142, g22);
not(t_143, f40);
or(t48, t_142, t_143);
not(u48, h38);
not(v48, i38);
buf(w48, j38);
not(x48, l38);
not(t_144, i22);
not(t_145, p40);
or(y48, t_144, t_145);
not(t_146, p38);
not(t_147, n38);
or(z48, t_146, t_147);
not(a49, n38);
not(b49, o38);
not(t_148, k22);
not(t_149, o40);
or(c49, t_148, t_149);
not(t_150, v38);
not(t_151, c33);
or(d49, t_150, t_151);
or(e49, a43, f18);
not(t_152, f18);
not(t_153, z42);
and(f49, t_152, t_153);
or(g49, y42, f18);
or(h49, b43, g18);
not(i49, r38);
not(j49, s38);
and(k49, x38, d33);
and(l49, w38, e33);
not(m49, t38);
and(n49, w38, e33);
and(o49, w38, e33);
not(p49, u38);
not(t_154, q38);
not(t_155, f33);
or(q49, t_154, t_155);
buf(r49, w38);
buf(s49, w38);
not(t49, x38);
not(u49, b39);
not(v49, c39);
not(t_156, t22);
not(t_157, x45);
or(w49, t_156, t_157);
not(t_158, u22);
not(t_159, y45);
or(x49, t_158, t_159);
not(t_160, v22);
not(t_161, h45);
or(y49, t_160, t_161);
not(t_162, w22);
not(t_163, i45);
or(z49, t_162, t_163);
not(a50, g39);
not(b50, h39);
not(t_164, y22);
not(t_165, n45);
or(c50, t_164, t_165);
not(d50, l39);
not(e50, m39);
not(t_166, a23);
not(t_167, o45);
or(f50, t_166, t_167);
buf(g50, n39);
not(h50, p39);
not(t_168, b23);
not(t_169, r45);
or(i50, t_168, t_169);
not(t_170, t39);
not(t_171, r39);
or(j50, t_170, t_171);
not(k50, r39);
not(l50, s39);
not(t_172, d23);
not(t_173, s45);
or(m50, t_172, t_173);
not(t_174, u39);
not(t_175, b40);
or(n50, t_174, t_175);
not(o50, v39);
not(p50, w39);
not(q50, x39);
not(r50, y39);
not(s50, z39);
not(t50, a40);
not(u50, b40);
not(v50, c40);
not(t_176, d40);
not(t_177, n40);
or(w50, t_176, t_177);
not(x50, e40);
not(y50, f40);
not(z50, g40);
not(a51, h40);
not(b51, i40);
not(c51, j40);
not(d51, k40);
not(e51, l40);
not(f51, m40);
not(g51, n40);
not(h51, o40);
not(i51, p40);
buf(j51, q40);
and(k51, l42, q40);
buf(l51, q40);
buf(m51, r40);
buf(n51, r40);
buf(o51, r40);
buf(p51, s40);
buf(q51, s40);
buf(r51, s40);
and(s51, k42, t40);
buf(t51, t40);
buf(u51, t40);
buf(v51, u40);
buf(w51, u40);
buf(x51, u40);
and(y51, j42, v40);
buf(z51, v40);
buf(a52, v40);
buf(b52, w40);
buf(c52, w40);
buf(d52, w40);
and(e52, p41, x40);
buf(f52, x40);
buf(g52, x40);
and(h52, t41, y40);
buf(i52, y40);
buf(j52, y40);
buf(k52, z40);
buf(l52, z40);
buf(m52, z40);
not(n52, a41);
not(o52, b41);
not(t_178, f29);
not(t_179, l45);
or(p52, t_178, t_179);
not(t_180, g29);
not(t_181, m45);
or(q52, t_180, t_181);
not(r52, f41);
not(s52, g41);
buf(t52, h41);
and(u52, x41, h41);
buf(v52, h41);
buf(w52, i41);
buf(x52, i41);
buf(y52, i41);
buf(z52, j41);
buf(a53, j41);
buf(b53, j41);
buf(c53, k41);
and(d53, i42, k41);
buf(e53, k41);
buf(f53, l41);
buf(g53, l41);
buf(h53, l41);
and(i53, s41, m41);
buf(j53, m41);
buf(k53, m41);
buf(l53, n41);
buf(m53, n41);
buf(n53, n41);
buf(o53, o41);
and(p53, g42, o41);
buf(q53, o41);
buf(r53, p41);
buf(s53, p41);
buf(t53, q41);
buf(u53, q41);
buf(v53, r41);
buf(w53, r41);
buf(x53, s41);
buf(y53, s41);
buf(z53, t41);
buf(a54, t41);
buf(b54, u41);
buf(c54, u41);
buf(d54, v41);
buf(e54, v41);
buf(f54, w41);
buf(g54, w41);
buf(h54, x41);
buf(i54, x41);
not(j54, y41);
not(k54, z41);
buf(l54, a42);
buf(m54, a42);
buf(n54, a42);
and(o54, d42, a35);
not(p54, b42);
not(q54, c42);
buf(r54, d42);
buf(s54, d42);
buf(t54, e42);
buf(u54, e42);
buf(v54, f42);
buf(w54, f42);
buf(x54, g42);
buf(y54, g42);
not(z54, h42);
buf(a55, i42);
buf(b55, i42);
buf(c55, j42);
buf(d55, j42);
buf(e55, k42);
buf(f55, k42);
buf(g55, l42);
buf(h55, l42);
buf(i55, m42);
buf(j55, m42);
buf(k55, m42);
and(l55, e42, b35);
not(m55, n42);
not(n55, o42);
and(o55, q41, c35);
not(p55, p42);
not(q55, q42);
buf(r55, r42);
buf(s55, r42);
buf(t55, r42);
not(t_182, s42);
not(t_183, u42);
or(u55, t_182, t_183);
not(v55, t42);
not(w55, u42);
buf(x55, v42);
and(y55, s36, z30);
not(t_184, f35);
not(t_185, w42);
or(z55, t_184, t_185);
not(t_186, i35);
not(t_187, r38);
or(a56, t_186, t_187);
not(t_188, c31);
not(t_189, s38);
or(b56, t_188, t_189);
and(c56, r41, l35);
not(d56, c43);
not(e56, d43);
buf(f56, e43);
buf(g56, e43);
buf(h56, e43);
buf(i56, f43);
buf(j56, f43);
buf(k56, f43);
and(l56, f42, m35);
not(m56, g43);
not(n56, h43);
buf(o56, i43);
buf(p56, i43);
buf(q56, i43);
and(r56, w41, n35);
not(s56, j43);
not(t56, k43);
buf(u56, l43);
buf(v56, l43);
buf(w56, l43);
not(x56, m43);
and(y56, u41, o35);
not(z56, n43);
buf(a57, o43);
buf(b57, o43);
buf(c57, o43);
and(d57, v41, p35);
not(e57, p43);
not(f57, q43);
and(g57, q35, u43);
not(h57, r43);
not(i57, s43);
not(j57, t43);
buf(k57, u43);
and(l57, v42, s15);
not(m57, v43);
not(n57, w43);
not(o57, x43);
not(p57, y43);
not(q57, z43);
not(r57, a44);
not(s57, b44);
not(t57, c44);
not(u57, d44);
not(t_190, f44);
not(t_191, x35);
or(v57, t_190, t_191);
not(t_192, e44);
not(t_193, y35);
or(w57, t_192, t_193);
not(x57, g44);
not(y57, h44);
not(z57, i44);
not(a58, j44);
not(b58, k44);
not(c58, l44);
not(d58, m44);
not(e58, n44);
not(f58, o44);
not(g58, p44);
not(h58, q44);
not(i58, r44);
not(j58, s44);
not(k58, t44);
not(l58, u44);
not(m58, v44);
not(n58, w44);
not(o58, x44);
not(p58, y44);
not(q58, z44);
not(r58, a45);
not(s58, b45);
not(t58, c45);
not(u58, d45);
not(v58, e45);
not(w58, f45);
not(x58, g45);
not(y58, h45);
not(z58, i45);
not(a59, j45);
not(b59, k45);
not(c59, l45);
not(d59, m45);
not(e59, n45);
not(f59, o45);
not(g59, p45);
not(h59, q45);
not(i59, r45);
not(j59, s45);
not(k59, t45);
not(t_194, v45);
not(t_195, p36);
or(l59, t_194, t_195);
not(t_196, u45);
not(t_197, q36);
or(m59, t_196, t_197);
not(n59, w45);
not(o59, x45);
not(p59, y45);
and(q59, z55, s36);
not(t_198, c20);
not(t_199, l54);
or(r59, t_198, t_199);
not(t_200, d20);
not(t_201, n54);
or(s59, t_200, t_201);
not(t_202, e20);
not(t_203, i55);
or(t59, t_202, t_203);
not(t_204, f20);
not(t_205, k55);
or(u59, t_204, t_205);
not(t_206, g20);
not(t_207, k56);
or(v59, t_206, t_207);
not(t_208, h20);
not(t_209, j56);
or(w59, t_208, t_209);
buf(x59, f46);
buf(y59, g46);
not(z59, h46);
not(t_210, i20);
not(t_211, g56);
or(a60, t_210, t_211);
not(t_212, j20);
not(t_213, h56);
or(b60, t_212, t_213);
not(c60, i46);
not(t_214, k20);
not(t_215, t55);
or(d60, t_214, t_215);
not(t_216, l20);
not(t_217, r55);
or(e60, t_216, t_217);
not(t_218, m20);
not(t_219, c52);
or(f60, t_218, t_219);
not(t_220, n20);
not(t_221, d52);
or(g60, t_220, t_221);
not(t_222, o20);
not(t_223, m53);
or(h60, t_222, t_223);
not(t_224, p20);
not(t_225, n53);
or(i60, t_224, t_225);
not(t_226, q20);
not(t_227, g53);
or(j60, t_226, t_227);
not(t_228, r20);
not(t_229, h53);
or(k60, t_228, t_229);
buf(l60, s46);
not(t_230, s20);
not(t_231, l52);
or(m60, t_230, t_231);
not(n60, t46);
not(t_232, t20);
not(t_233, m52);
or(o60, t_232, t_233);
not(t_234, u20);
not(t_235, a53);
or(p60, t_234, t_235);
not(t_236, v20);
not(t_237, b53);
or(q60, t_236, t_237);
not(t_238, w20);
not(t_239, v51);
or(r60, t_238, t_239);
not(t_240, x20);
not(t_241, w51);
or(s60, t_240, t_241);
not(t_242, y20);
not(t_243, q51);
or(t60, t_242, t_243);
not(t_244, z20);
not(t_245, r51);
or(u60, t_244, t_245);
buf(v60, a47);
buf(w60, b47);
not(x60, c47);
not(t_246, a21);
not(t_247, n51);
or(y60, t_246, t_247);
not(t_248, b21);
not(t_249, m51);
or(z60, t_248, t_249);
not(a61, d47);
not(t_250, c21);
not(t_251, y52);
or(b61, t_250, t_251);
not(t_252, d21);
not(t_253, x52);
or(c61, t_252, t_253);
not(t_254, e21);
not(t_255, b57);
or(d61, t_254, t_255);
not(t_256, f21);
not(t_257, a57);
or(e61, t_256, t_257);
not(t_258, g21);
not(t_259, w56);
or(f61, t_258, t_259);
not(t_260, h21);
not(t_261, v56);
or(g61, t_260, t_261);
not(t_262, i21);
not(t_263, p56);
or(h61, t_262, t_263);
not(t_264, j21);
not(t_265, o56);
or(i61, t_264, t_265);
not(t_266, q47);
not(t_267, u36);
or(j61, t_266, t_267);
not(t_268, a58);
not(t_269, v36);
or(k61, t_268, t_269);
not(t_270, t58);
not(t_271, n17);
or(l61, t_270, t_271);
not(t_272, u58);
not(t_273, o17);
or(m61, t_272, t_273);
not(t_274, m47);
not(t_275, z36);
or(n61, t_274, t_275);
not(t_276, b58);
not(t_277, a37);
or(o61, t_276, t_277);
not(t_278, v58);
not(t_279, p17);
or(p61, t_278, t_279);
not(t_280, w58);
not(t_281, q17);
or(q61, t_280, t_281);
not(t_282, e58);
not(t_283, g37);
or(r61, t_282, t_283);
not(t_284, e48);
not(t_285, h37);
or(s61, t_284, t_285);
not(t_286, l58);
not(t_287, r17);
or(t61, t_286, t_287);
not(t_288, k58);
not(t_289, s17);
or(u61, t_288, t_289);
not(v61, y47);
not(w61, z47);
not(t_290, n58);
not(t_291, t17);
or(x61, t_290, t_291);
not(t_292, m58);
not(t_293, u17);
or(y61, t_292, t_293);
not(t_294, v47);
not(t_295, n37);
or(z61, t_294, t_295);
not(t_296, f58);
not(t_297, o37);
or(a62, t_296, t_297);
not(t_298, n48);
not(t_299, q37);
or(b62, t_298, t_299);
not(t_300, i58);
not(t_301, r37);
or(c62, t_300, t_301);
not(t_302, r58);
not(t_303, v17);
or(d62, t_302, t_303);
not(t_304, q58);
not(t_305, w17);
or(e62, t_304, t_305);
not(t_306, f51);
not(t_307, x17);
or(f62, t_306, t_307);
not(t_308, e51);
not(t_309, y17);
or(g62, t_308, t_309);
not(t_310, s50);
not(t_311, x37);
or(h62, t_310, t_311);
not(t_312, g48);
not(t_313, y37);
or(i62, t_312, t_313);
not(t_314, v48);
not(t_315, c38);
or(j62, t_314, t_315);
not(t_316, r50);
not(t_317, d38);
or(k62, t_316, t_317);
not(t_318, c51);
not(t_319, z17);
or(l62, t_318, t_319);
not(t_320, b51);
not(t_321, a18);
or(m62, t_320, t_321);
not(t_322, z50);
not(t_323, b18);
or(n62, t_322, t_323);
not(t_324, y50);
not(t_325, c18);
or(o62, t_324, t_325);
not(t_326, o50);
not(t_327, h38);
or(p62, t_326, t_327);
not(t_328, o48);
not(t_329, i38);
or(q62, t_328, t_329);
not(r62, w48);
not(t_330, i51);
not(t_331, d18);
or(s62, t_330, t_331);
not(t_332, v50);
not(t_333, o38);
or(t62, t_332, t_333);
not(t_334, h51);
not(t_335, e18);
or(u62, t_334, t_335);
not(t_336, a49);
not(t_337, b33);
or(v62, t_336, t_337);
not(t_338, d49);
not(t_339, q49);
or(w62, t_338, t_339);
or(x62, l49, e49);
not(y62, e49);
not(z62, f49);
not(a63, g49);
or(b63, o49, x42, f18);
not(c63, h49);
not(d63, k49);
not(e63, n49);
not(f63, r49);
not(g63, s49);
not(t_340, b50);
not(t_341, b39);
or(h63, t_340, t_341);
not(t_342, y57);
not(t_343, c39);
or(i63, t_342, t_343);
not(t_344, o59);
not(t_345, k18);
or(j63, t_344, t_345);
not(t_346, p59);
not(t_347, l18);
or(k63, t_346, t_347);
not(t_348, y58);
not(t_349, m18);
or(l63, t_348, t_349);
not(t_350, z58);
not(t_351, n18);
or(m63, t_350, t_351);
not(t_352, o57);
not(t_353, g39);
or(n63, t_352, t_353);
not(t_354, u49);
not(t_355, h39);
or(o63, t_354, t_355);
not(t_356, e59);
not(t_357, o18);
or(p63, t_356, t_357);
not(t_358, s57);
not(t_359, l39);
or(q63, t_358, t_359);
not(t_360, r52);
not(t_361, m39);
or(r63, t_360, t_361);
not(t_362, f59);
not(t_363, p18);
or(s63, t_362, t_363);
not(t63, g50);
not(t_364, i59);
not(t_365, q18);
or(u63, t_364, t_365);
not(t_366, u57);
not(t_367, s39);
or(v63, t_366, t_367);
not(t_368, j59);
not(t_369, r18);
or(w63, t_368, t_369);
not(t_370, k50);
not(t_371, k33);
or(x63, t_370, t_371);
not(t_372, u50);
not(t_373, p34);
or(y63, t_372, t_373);
not(t_374, u48);
not(t_375, v39);
or(z63, t_374, t_375);
not(t_376, q50);
not(t_377, w39);
or(a64, t_376, t_377);
not(t_378, p50);
not(t_379, x39);
or(b64, t_378, t_379);
not(t_380, p48);
not(t_381, y39);
or(c64, t_380, t_381);
not(t_382, m48);
not(t_383, z39);
or(d64, t_382, t_383);
not(t_384, h58);
not(t_385, a40);
or(e64, t_384, t_385);
not(t_386, b49);
not(t_387, c40);
or(f64, t_386, t_387);
not(t_388, g51);
not(t_389, u34);
or(g64, t_388, t_389);
not(t_390, a51);
not(t_391, e40);
or(h64, t_390, t_391);
not(t_392, x50);
not(t_393, h40);
or(i64, t_392, t_393);
not(t_394, p58);
not(t_395, k40);
or(j64, t_394, t_395);
not(k64, j51);
not(l64, l51);
not(m64, m51);
not(n64, n51);
not(o64, o51);
not(p64, p51);
not(q64, q51);
not(r64, r51);
not(s64, t51);
not(t64, u51);
not(u64, v51);
not(v64, w51);
not(w64, x51);
not(x64, z51);
not(y64, a52);
not(z64, b52);
not(a65, c52);
not(b65, d52);
not(c65, f52);
not(t_396, q55);
not(t_397, g52);
or(d65, t_396, t_397);
not(e65, g52);
not(f65, i52);
not(t_398, n52);
not(t_399, j52);
or(g65, t_398, t_399);
not(h65, j52);
not(t_400, o52);
not(t_401, k52);
or(i65, t_400, t_401);
not(j65, k52);
not(k65, l52);
not(l65, m52);
not(t_402, c59);
not(t_403, n24);
or(m65, t_402, t_403);
not(t_404, d59);
not(t_405, o24);
or(n65, t_404, t_405);
not(t_406, e50);
not(t_407, f41);
or(o65, t_406, t_407);
not(t_408, q57);
not(t_409, g41);
or(p65, t_408, t_409);
not(q65, t52);
not(t_410, f57);
not(t_411, v52);
or(r65, t_410, t_411);
not(s65, v52);
not(t65, w52);
not(u65, x52);
not(v65, y52);
not(w65, z52);
not(x65, a53);
not(y65, b53);
not(z65, c53);
not(a66, e53);
not(b66, f53);
not(c66, g53);
not(d66, h53);
not(e66, j53);
not(f66, k53);
not(g66, l53);
not(h66, m53);
not(i66, n53);
not(j66, o53);
not(k66, q53);
not(l66, r53);
not(m66, s53);
not(t_412, p55);
not(t_413, t53);
or(n66, t_412, t_413);
not(o66, t53);
not(p66, u53);
not(t_414, d56);
not(t_415, v53);
or(q66, t_414, t_415);
not(r66, v53);
not(s66, w53);
not(t66, x53);
not(u66, y53);
not(v66, z53);
not(t_416, z54);
not(t_417, a54);
or(w66, t_416, t_417);
not(x66, a54);
not(y66, b54);
not(t_418, x56);
not(t_419, c54);
or(z66, t_418, t_419);
not(a67, c54);
not(t_420, e57);
not(t_421, d54);
or(b67, t_420, t_421);
not(c67, d54);
not(d67, e54);
not(t_422, s56);
not(t_423, f54);
or(e67, t_422, t_423);
not(f67, f54);
not(g67, g54);
not(h67, h54);
not(i67, i54);
not(t_424, k54);
not(t_425, y41);
or(j67, t_424, t_425);
not(t_426, j54);
not(t_427, z41);
or(k67, t_426, t_427);
not(l67, l54);
not(m67, m54);
not(n67, n54);
not(t_428, n55);
not(t_429, b42);
or(o67, t_428, t_429);
not(t_430, q54);
not(t_431, r54);
or(p67, t_430, t_431);
not(q67, r54);
not(r67, s54);
not(t_432, m55);
not(t_433, t54);
or(s67, t_432, t_433);
not(t67, t54);
not(u67, u54);
not(t_434, m56);
not(t_435, v54);
or(v67, t_434, t_435);
not(w67, v54);
not(x67, w54);
not(y67, x54);
not(z67, y54);
not(a68, a55);
not(b68, b55);
not(c68, c55);
not(d68, d55);
not(e68, e55);
not(f68, f55);
not(g68, g55);
not(h68, h55);
not(i68, i55);
not(j68, j55);
not(k68, k55);
not(t_436, p54);
not(t_437, o42);
or(l68, t_436, t_437);
not(m68, r55);
not(n68, s55);
not(o68, t55);
not(t_438, w55);
not(t_439, d35);
or(p68, t_438, t_439);
not(t_440, v55);
not(t_441, x55);
or(q68, t_440, t_441);
not(r68, x55);
or(s68, y55, w24);
not(t_442, i49);
not(t_443, b31);
or(t68, t_442, t_443);
not(t_444, j49);
not(t_445, a25);
or(u68, t_444, t_445);
not(t_446, n56);
not(t_447, d43);
or(v68, t_446, t_447);
not(w68, f56);
not(x68, g56);
not(y68, h56);
not(z68, i56);
not(a69, j56);
not(b69, k56);
not(t_448, e56);
not(t_449, h43);
or(c69, t_448, t_449);
not(d69, o56);
not(e69, p56);
not(f69, q56);
not(t_450, z56);
not(t_451, k43);
or(g69, t_450, t_451);
not(h69, u56);
not(i69, v56);
not(j69, w56);
not(t_452, t56);
not(t_453, n43);
or(k69, t_452, t_453);
not(l69, a57);
not(m69, b57);
not(n69, c57);
not(t_454, h57);
not(t_455, k57);
or(o69, t_454, t_455);
and(p69, r35, l57);
and(q69, r35, l57);
not(t_456, r35);
not(t_457, l57);
and(r69, t_456, t_457);
not(s69, k57);
buf(t69, l57);
buf(u69, l57);
not(t_458, t57);
not(t_459, v43);
or(v69, t_458, t_459);
not(t_460, x57);
not(t_461, w43);
or(w69, t_460, t_461);
not(t_462, a50);
not(t_463, x43);
or(x69, t_462, t_463);
not(t_464, r57);
not(t_465, y43);
or(y69, t_464, t_465);
not(t_466, s52);
not(t_467, z43);
or(z69, t_466, t_467);
not(t_468, p57);
not(t_469, a44);
or(a70, t_468, t_469);
not(t_470, d50);
not(t_471, b44);
or(b70, t_470, t_471);
not(t_472, m57);
not(t_473, c44);
or(c70, t_472, t_473);
not(t_474, l50);
not(t_475, d44);
or(d70, t_474, t_475);
not(t_476, v57);
not(t_477, w57);
or(e70, t_476, t_477);
not(t_478, n57);
not(t_479, g44);
or(f70, t_478, t_479);
not(t_480, v49);
not(t_481, h44);
or(g70, t_480, t_481);
not(t_482, c58);
not(t_483, i44);
or(h70, t_482, t_483);
not(t_484, n47);
not(t_485, j44);
or(i70, t_484, t_485);
not(t_486, r47);
not(t_487, k44);
or(j70, t_486, t_487);
not(t_488, z57);
not(t_489, l44);
or(k70, t_488, t_489);
not(t_490, g58);
not(t_491, m44);
or(l70, t_490, t_491);
not(t_492, u47);
not(t_493, n44);
or(m70, t_492, t_493);
not(t_494, f48);
not(t_495, o44);
or(n70, t_494, t_495);
not(t_496, d58);
not(t_497, p44);
or(o70, t_496, t_497);
not(t_498, t50);
not(t_499, q44);
or(p70, t_498, t_499);
not(t_500, h48);
not(t_501, r44);
or(q70, t_500, t_501);
not(t_502, o58);
not(t_503, s44);
or(r70, t_502, t_503);
not(t_504, j58);
not(t_505, x44);
or(s70, t_504, t_505);
not(t_506, d51);
not(t_507, y44);
or(t70, t_506, t_507);
not(t_508, x58);
not(t_509, b45);
or(u70, t_508, t_509);
not(t_510, s58);
not(t_511, g45);
or(v70, t_510, t_511);
not(t_512, n59);
not(t_513, j45);
or(w70, t_512, t_513);
not(t_514, g59);
not(t_515, k45);
or(x70, t_514, t_515);
not(t_516, b59);
not(t_517, p45);
or(y70, t_516, t_517);
not(t_518, k59);
not(t_519, q45);
or(z70, t_518, t_519);
not(t_520, h59);
not(t_521, t45);
or(a71, t_520, t_521);
not(t_522, l59);
not(t_523, m59);
or(b71, t_522, t_523);
not(t_524, a59);
not(t_525, w45);
or(c71, t_524, t_525);
not(d71, q59);
not(t_526, l67);
not(t_527, f16);
or(e71, t_526, t_527);
not(t_528, n67);
not(t_529, g16);
or(f71, t_528, t_529);
not(t_530, i68);
not(t_531, h16);
or(g71, t_530, t_531);
not(t_532, k68);
not(t_533, i16);
or(h71, t_532, t_533);
not(t_534, b69);
not(t_535, j16);
or(i71, t_534, t_535);
not(t_536, a69);
not(t_537, k16);
or(j71, t_536, t_537);
not(k71, x59);
not(l71, y59);
not(t_538, x68);
not(t_539, l16);
or(m71, t_538, t_539);
not(t_540, y68);
not(t_541, m16);
or(n71, t_540, t_541);
not(t_542, o68);
not(t_543, n16);
or(o71, t_542, t_543);
not(t_544, m68);
not(t_545, o16);
or(p71, t_544, t_545);
not(t_546, a65);
not(t_547, p16);
or(q71, t_546, t_547);
not(t_548, b65);
not(t_549, q16);
or(r71, t_548, t_549);
not(t_550, h66);
not(t_551, r16);
or(s71, t_550, t_551);
not(t_552, i66);
not(t_553, s16);
or(t71, t_552, t_553);
not(t_554, c66);
not(t_555, t16);
or(u71, t_554, t_555);
not(t_556, d66);
not(t_557, u16);
or(v71, t_556, t_557);
not(w71, l60);
not(t_558, k65);
not(t_559, v16);
or(x71, t_558, t_559);
not(t_560, l65);
not(t_561, w16);
or(y71, t_560, t_561);
not(t_562, x65);
not(t_563, x16);
or(z71, t_562, t_563);
not(t_564, y65);
not(t_565, y16);
or(a72, t_564, t_565);
not(t_566, u64);
not(t_567, z16);
or(b72, t_566, t_567);
not(t_568, v64);
not(t_569, a17);
or(c72, t_568, t_569);
not(t_570, q64);
not(t_571, b17);
or(d72, t_570, t_571);
not(t_572, r64);
not(t_573, c17);
or(e72, t_572, t_573);
not(f72, v60);
not(g72, w60);
not(t_574, n64);
not(t_575, d17);
or(h72, t_574, t_575);
not(t_576, m64);
not(t_577, e17);
or(i72, t_576, t_577);
not(t_578, v65);
not(t_579, f17);
or(j72, t_578, t_579);
not(t_580, u65);
not(t_581, g17);
or(k72, t_580, t_581);
not(t_582, m69);
not(t_583, h17);
or(l72, t_582, t_583);
not(t_584, l69);
not(t_585, i17);
or(m72, t_584, t_585);
not(t_586, j69);
not(t_587, j17);
or(n72, t_586, t_587);
not(t_588, i69);
not(t_589, k17);
or(o72, t_588, t_589);
not(t_590, e69);
not(t_591, l17);
or(p72, t_590, t_591);
not(t_592, d69);
not(t_593, m17);
or(q72, t_592, t_593);
not(t_594, j61);
not(t_595, n61);
or(r72, t_594, t_595);
not(t_596, k61);
not(t_597, i70);
or(s72, t_596, t_597);
not(t_598, l61);
not(t_599, o47);
or(t72, t_598, t_599);
not(t_600, m61);
not(t_601, p47);
or(u72, t_600, t_601);
not(t_602, o61);
not(t_603, j70);
or(v72, t_602, t_603);
not(t_604, p61);
not(t_605, s47);
or(w72, t_604, t_605);
not(t_606, q61);
not(t_607, t47);
or(x72, t_606, t_607);
not(t_608, r61);
not(t_609, m70);
or(y72, t_608, t_609);
not(t_610, s61);
not(t_611, z61);
or(z72, t_610, t_611);
not(t_612, t61);
not(t_613, w47);
or(a73, t_612, t_613);
not(t_614, u61);
not(t_615, x47);
or(b73, t_614, t_615);
not(t_616, x61);
not(t_617, a48);
or(c73, t_616, t_617);
not(t_618, y61);
not(t_619, d48);
or(d73, t_618, t_619);
not(t_620, a62);
not(t_621, n70);
or(e73, t_620, t_621);
not(t_622, b62);
not(t_623, i62);
or(f73, t_622, t_623);
not(t_624, c62);
not(t_625, q70);
or(g73, t_624, t_625);
not(t_626, d62);
not(t_627, i48);
or(h73, t_626, t_627);
not(t_628, e62);
not(t_629, j48);
or(i73, t_628, t_629);
not(t_630, f62);
not(t_631, k48);
or(j73, t_630, t_631);
not(t_632, g62);
not(t_633, l48);
or(k73, t_632, t_633);
not(t_634, h62);
not(t_635, d64);
or(l73, t_634, t_635);
not(t_636, j62);
not(t_637, q62);
or(m73, t_636, t_637);
not(t_638, k62);
not(t_639, c64);
or(n73, t_638, t_639);
not(t_640, l62);
not(t_641, q48);
or(o73, t_640, t_641);
not(t_642, m62);
not(t_643, r48);
or(p73, t_642, t_643);
not(t_644, n62);
not(t_645, s48);
or(q73, t_644, t_645);
not(t_646, o62);
not(t_647, t48);
or(r73, t_646, t_647);
not(t_648, p62);
not(t_649, z63);
or(s73, t_648, t_649);
not(t_650, s62);
not(t_651, y48);
or(t73, t_650, t_651);
not(t_652, z48);
not(t_653, v62);
or(u73, t_652, t_653);
not(t_654, t62);
not(t_655, f64);
or(v73, t_654, t_655);
not(t_656, u62);
not(t_657, c49);
or(w73, t_656, t_657);
not(x73, w62);
not(y73, x62);
not(z73, y62);
not(t_658, e63);
not(t_659, a63);
or(a74, t_658, t_659);
not(b74, b63);
not(t_660, d63);
not(t_661, c63);
or(c74, t_660, t_661);
not(t_662, h63);
not(t_663, o63);
or(d74, t_662, t_663);
not(t_664, i63);
not(t_665, g70);
or(e74, t_664, t_665);
not(t_666, j63);
not(t_667, w49);
or(f74, t_666, t_667);
not(t_668, k63);
not(t_669, x49);
or(g74, t_668, t_669);
not(t_670, l63);
not(t_671, y49);
or(h74, t_670, t_671);
not(t_672, m63);
not(t_673, z49);
or(i74, t_672, t_673);
not(t_674, n63);
not(t_675, x69);
or(j74, t_674, t_675);
not(t_676, p63);
not(t_677, c50);
or(k74, t_676, t_677);
not(t_678, q63);
not(t_679, b70);
or(l74, t_678, t_679);
not(t_680, o65);
not(t_681, r63);
or(m74, t_680, t_681);
not(t_682, s63);
not(t_683, f50);
or(n74, t_682, t_683);
not(t_684, u63);
not(t_685, i50);
or(o74, t_684, t_685);
not(t_686, j50);
not(t_687, x63);
or(p74, t_686, t_687);
not(t_688, v63);
not(t_689, d70);
or(q74, t_688, t_689);
not(t_690, w63);
not(t_691, m50);
or(r74, t_690, t_691);
not(t_692, n50);
not(t_693, y63);
or(s74, t_692, t_693);
not(t_694, b64);
not(t_695, a64);
or(t74, t_694, t_695);
not(t_696, p70);
not(t_697, e64);
or(u74, t_696, t_697);
not(t_698, w50);
not(t_699, g64);
or(v74, t_698, t_699);
not(t_700, i64);
not(t_701, h64);
or(w74, t_700, t_701);
not(t_702, t70);
not(t_703, j64);
or(x74, t_702, t_703);
not(t_704, t64);
not(t_705, j51);
or(y74, t_704, t_705);
not(t_706, h68);
not(t_707, l51);
or(z74, t_706, t_707);
not(t_708, p64);
not(t_709, o51);
or(a75, t_708, t_709);
not(t_710, o64);
not(t_711, p51);
or(b75, t_710, t_711);
not(t_712, f68);
not(t_713, t51);
or(c75, t_712, t_713);
not(t_714, k64);
not(t_715, u51);
or(d75, t_714, t_715);
not(t_716, w65);
not(t_717, x51);
or(e75, t_716, t_717);
not(t_718, c68);
not(t_719, z51);
or(f75, t_718, t_719);
not(t_720, a66);
not(t_721, a52);
or(g75, t_720, t_721);
not(t_722, n68);
not(t_723, b52);
or(h75, t_722, t_723);
not(t_724, l66);
not(t_725, f52);
or(i75, t_724, t_725);
not(t_726, v66);
not(t_727, i52);
or(j75, t_726, t_727);
not(t_728, h65);
not(t_729, a41);
or(k75, t_728, t_729);
not(t_730, j65);
not(t_731, b41);
or(l75, t_730, t_731);
not(t_732, m65);
not(t_733, p52);
or(m75, t_732, t_733);
not(t_734, n65);
not(t_735, q52);
or(n75, t_734, t_735);
not(t_736, p65);
not(t_737, z69);
or(o75, t_736, t_737);
not(t_738, i67);
not(t_739, t52);
or(p75, t_738, t_739);
not(t_740, n69);
not(t_741, w52);
or(q75, t_740, t_741);
not(t_742, w64);
not(t_743, z52);
or(r75, t_742, t_743);
not(t_744, b68);
not(t_745, c53);
or(s75, t_744, t_745);
not(t_746, y64);
not(t_747, e53);
or(t75, t_746, t_747);
not(t_748, g66);
not(t_749, f53);
or(u75, t_748, t_749);
not(t_750, t66);
not(t_751, j53);
or(v75, t_750, t_751);
not(t_752, k66);
not(t_753, k53);
or(w75, t_752, t_753);
not(t_754, b66);
not(t_755, l53);
or(x75, t_754, t_755);
not(t_756, y67);
not(t_757, o53);
or(y75, t_756, t_757);
not(t_758, f66);
not(t_759, q53);
or(z75, t_758, t_759);
not(t_760, c65);
not(t_761, r53);
or(a76, t_760, t_761);
not(t_762, p66);
not(t_763, s53);
or(b76, t_762, t_763);
not(t_764, m66);
not(t_765, u53);
or(c76, t_764, t_765);
not(t_766, x67);
not(t_767, w53);
or(d76, t_766, t_767);
not(t_768, e66);
not(t_769, x53);
or(e76, t_768, t_769);
not(t_770, z67);
not(t_771, y53);
or(f76, t_770, t_771);
not(t_772, f65);
not(t_773, z53);
or(g76, t_772, t_773);
not(t_774, g67);
not(t_775, b54);
or(h76, t_774, t_775);
not(t_776, h67);
not(t_777, e54);
or(i76, t_776, t_777);
not(t_778, y66);
not(t_779, g54);
or(j76, t_778, t_779);
not(t_780, d67);
not(t_781, h54);
or(k76, t_780, t_781);
not(t_782, q65);
not(t_783, i54);
or(l76, t_782, t_783);
not(t_784, j67);
not(t_785, k67);
or(m76, t_784, t_785);
not(t_786, j68);
not(t_787, m54);
or(n76, t_786, t_787);
not(t_788, o67);
not(t_789, l68);
or(o76, t_788, t_789);
not(t_790, q67);
not(t_791, c42);
or(p76, t_790, t_791);
not(t_792, u67);
not(t_793, s54);
or(q76, t_792, t_793);
not(t_794, r67);
not(t_795, u54);
or(r76, t_794, t_795);
not(t_796, s66);
not(t_797, w54);
or(s76, t_796, t_797);
not(t_798, j66);
not(t_799, x54);
or(t76, t_798, t_799);
not(t_800, u66);
not(t_801, y54);
or(u76, t_800, t_801);
not(t_802, x66);
not(t_803, h42);
or(v76, t_802, t_803);
not(t_804, d68);
not(t_805, a55);
or(w76, t_804, t_805);
not(t_806, z65);
not(t_807, b55);
or(x76, t_806, t_807);
not(t_808, x64);
not(t_809, c55);
or(y76, t_808, t_809);
not(t_810, a68);
not(t_811, d55);
or(z76, t_810, t_811);
not(t_812, g68);
not(t_813, e55);
or(a77, t_812, t_813);
not(t_814, s64);
not(t_815, f55);
or(b77, t_814, t_815);
not(t_816, e68);
not(t_817, g55);
or(c77, t_816, t_817);
not(t_818, l64);
not(t_819, h55);
or(d77, t_818, t_819);
not(t_820, m67);
not(t_821, j55);
or(e77, t_820, t_821);
not(t_822, t67);
not(t_823, n42);
or(f77, t_822, t_823);
not(t_824, o66);
not(t_825, p42);
or(g77, t_824, t_825);
not(t_826, e65);
not(t_827, q42);
or(h77, t_826, t_827);
not(t_828, z64);
not(t_829, s55);
or(i77, t_828, t_829);
not(t_830, u55);
not(t_831, p68);
or(j77, t_830, t_831);
not(t_832, r68);
not(t_833, t42);
or(k77, t_832, t_833);
not(l77, s68);
not(t_834, h35);
not(t_835, y62);
or(m77, t_834, t_835);
not(t_836, t68);
not(t_837, a56);
or(n77, t_836, t_837);
not(t_838, u68);
not(t_839, b56);
or(o77, t_838, t_839);
not(t_840, e31);
not(t_841, x62);
or(p77, t_840, t_841);
not(t_842, r66);
not(t_843, c43);
or(q77, t_842, t_843);
not(t_844, c69);
not(t_845, v68);
or(r77, t_844, t_845);
not(t_846, z68);
not(t_847, f56);
or(s77, t_846, t_847);
not(t_848, w68);
not(t_849, i56);
or(t77, t_848, t_849);
not(t_850, w67);
not(t_851, g43);
or(u77, t_850, t_851);
not(t_852, h69);
not(t_853, q56);
or(v77, t_852, t_853);
not(t_854, f67);
not(t_855, j43);
or(w77, t_854, t_855);
not(t_856, k69);
not(t_857, g69);
or(x77, t_856, t_857);
not(t_858, f69);
not(t_859, u56);
or(y77, t_858, t_859);
not(t_860, a67);
not(t_861, m43);
or(z77, t_860, t_861);
not(t_862, t65);
not(t_863, c57);
or(a78, t_862, t_863);
not(t_864, c67);
not(t_865, p43);
or(b78, t_864, t_865);
not(t_866, s65);
not(t_867, q43);
or(c78, t_866, t_867);
not(t_868, s69);
not(t_869, r43);
or(d78, t_868, t_869);
buf(e78, q69);
not(t_870, i57);
not(t_871, u69);
or(f78, t_870, t_871);
not(g78, r69);
not(t_872, j57);
not(t_873, t69);
or(h78, t_872, t_873);
not(i78, t69);
not(j78, u69);
not(t_874, c70);
not(t_875, v69);
or(k78, t_874, t_875);
not(t_876, f70);
not(t_877, w69);
or(l78, t_876, t_877);
not(t_878, y69);
not(t_879, a70);
or(m78, t_878, t_879);
not(n78, e70);
not(t_880, h70);
not(t_881, k70);
or(o78, t_880, t_881);
not(t_882, l70);
not(t_883, o70);
or(p78, t_882, t_883);
not(t_884, r70);
not(t_885, s70);
or(q78, t_884, t_885);
not(t_886, u70);
not(t_887, v70);
or(r78, t_886, t_887);
not(t_888, c71);
not(t_889, w70);
or(s78, t_888, t_889);
not(t_890, x70);
not(t_891, y70);
or(t78, t_890, t_891);
not(t_892, z70);
not(t_893, a71);
or(u78, t_892, t_893);
not(v78, b71);
not(t_894, d71);
not(t_895, l77);
or(w78, t_894, t_895);
not(t_896, e71);
not(t_897, r59);
or(x78, t_896, t_897);
not(t_898, f71);
not(t_899, s59);
or(y78, t_898, t_899);
not(t_900, g71);
not(t_901, t59);
or(z78, t_900, t_901);
not(t_902, h71);
not(t_903, u59);
or(a79, t_902, t_903);
not(t_904, i71);
not(t_905, v59);
or(b79, t_904, t_905);
not(t_906, j71);
not(t_907, w59);
or(c79, t_906, t_907);
not(t_908, m71);
not(t_909, a60);
or(d79, t_908, t_909);
not(t_910, n71);
not(t_911, b60);
or(e79, t_910, t_911);
not(t_912, o71);
not(t_913, d60);
or(f79, t_912, t_913);
not(t_914, p71);
not(t_915, e60);
or(g79, t_914, t_915);
not(t_916, q71);
not(t_917, f60);
or(h79, t_916, t_917);
not(t_918, r71);
not(t_919, g60);
or(i79, t_918, t_919);
not(t_920, s71);
not(t_921, h60);
or(j79, t_920, t_921);
not(t_922, t71);
not(t_923, i60);
or(k79, t_922, t_923);
not(t_924, u71);
not(t_925, j60);
or(l79, t_924, t_925);
not(t_926, v71);
not(t_927, k60);
or(m79, t_926, t_927);
not(t_928, x71);
not(t_929, m60);
or(n79, t_928, t_929);
not(t_930, y71);
not(t_931, o60);
or(o79, t_930, t_931);
not(t_932, z71);
not(t_933, p60);
or(p79, t_932, t_933);
not(t_934, a72);
not(t_935, q60);
or(q79, t_934, t_935);
not(t_936, b72);
not(t_937, r60);
or(r79, t_936, t_937);
not(t_938, c72);
not(t_939, s60);
or(s79, t_938, t_939);
not(t_940, d72);
not(t_941, t60);
or(t79, t_940, t_941);
not(t_942, e72);
not(t_943, u60);
or(u79, t_942, t_943);
not(t_944, h72);
not(t_945, y60);
or(v79, t_944, t_945);
not(t_946, i72);
not(t_947, z60);
or(w79, t_946, t_947);
not(t_948, j72);
not(t_949, b61);
or(x79, t_948, t_949);
not(t_950, k72);
not(t_951, c61);
or(y79, t_950, t_951);
not(t_952, l72);
not(t_953, d61);
or(z79, t_952, t_953);
not(t_954, m72);
not(t_955, e61);
or(a80, t_954, t_955);
not(t_956, n72);
not(t_957, f61);
or(b80, t_956, t_957);
not(t_958, o72);
not(t_959, g61);
or(c80, t_958, t_959);
not(t_960, p72);
not(t_961, h61);
or(d80, t_960, t_961);
not(t_962, q72);
not(t_963, i61);
or(e80, t_962, t_963);
not(f80, r72);
and(g80, e73, y72, v72, s72);
and(h80, d73, a73, x72, t72);
buf(i80, t72);
buf(j80, t72);
buf(k80, u72);
buf(l80, u72);
and(m80, w72, c73, b73, u72);
and(n80, s72, y36);
and(o80, u72, b37);
buf(p80, w72);
buf(q80, w72);
and(r80, c73, b73, w72);
and(s80, t72, c37);
buf(t80, x72);
and(u80, d73, a73, x72);
buf(v80, x72);
and(w80, x72, d37);
and(x80, x72, t72, d37);
and(y80, x72, d37);
and(z80, w72, u72, e37);
and(a81, w72, e37);
and(b81, w72, e37);
and(c81, v72, s72, f37);
not(d81, z72);
and(e81, d73, a73);
buf(f81, a73);
buf(g81, a73);
buf(h81, b73);
buf(i81, b73);
and(j81, c73, b73);
and(k81, a73, i37, x72);
and(l81, a73, t72, i37, x72);
and(m81, a73, i37, x72);
and(n81, a73, i37);
and(o81, b73, u72, j37, w72);
and(p81, j37, b73, w72);
and(q81, b73, j37, w72);
and(r81, b73, j37);
and(s81, b73, j37);
not(t81, c73);
buf(u81, d73);
buf(v81, d73);
and(w81, y72, s72, m37, v72);
buf(x81, f73);
buf(y81, f73);
and(z81, v73, s73, n73, l73, g73);
buf(a82, h73);
buf(b82, h73);
and(c82, t73, r73, o73, k73, h73);
and(d82, j73, w73, p73, i73, q73);
buf(e82, i73);
and(f82, h73, u37);
and(g82, i73, v37);
buf(h82, j73);
buf(i82, k73);
and(j82, t73, o73, k73, r73);
buf(k82, k73);
and(l82, g73, w37);
and(m82, k73, z37);
and(n82, k73, z37);
and(o82, k73, h73, z37);
and(p82, j73, a38);
and(q82, j73, i73, a38);
and(r82, l73, g73, b38);
not(s82, m73);
buf(t82, o73);
buf(u82, o73);
and(v82, t73, o73, r73);
buf(w82, p73);
and(x82, o73, e38, k73);
and(y82, o73, e38, k73);
and(z82, o73, h73, e38, k73);
and(a83, o73, e38);
and(b83, o73, e38);
and(c83, p73, f38, j73);
and(d83, p73, i73, f38, j73);
and(e83, f38, p73);
buf(f83, q73);
buf(g83, r73);
buf(h83, r73);
and(i83, t73, r73);
and(j83, n73, g73, g38, l73);
and(k83, r73, o73, j38, k73);
and(l83, r73, o73, h73, j38, k73);
and(m83, r73, o73, j38, k73);
and(n83, r73, o73, j38);
and(o83, r73, j38);
and(p83, r73, o73, j38);
and(q83, q73, p73, k38, j73);
and(r83, q73, p73, i73, k38, j73);
and(s83, q73, k38);
and(t83, q73, p73, k38);
buf(u83, t73);
buf(v83, t73);
and(w83, s73, n73, g73, m38, l73);
not(x83, u73);
buf(y83, w73);
buf(z83, d74);
buf(a84, d74);
and(b84, q74, l74, o75, j74, e74);
buf(c84, f74);
buf(d84, f74);
and(e84, o74, n74, m75, i74, f74);
and(f84, h74, r74, n75, g74, k74);
buf(g84, g74);
and(h84, f74, d39);
and(i84, g74, e39);
buf(j84, h74);
buf(k84, i74);
and(l84, o74, m75, i74, n74);
buf(m84, i74);
and(n84, e74, f39);
and(o84, m75, i39, i74);
and(p84, m75, i39, i74);
and(q84, m75, f74, i39, i74);
and(r84, m75, i39);
and(s84, m75, i39);
and(t84, n75, j39, h74);
and(u84, n75, g74, j39, h74);
and(v84, j39, n75);
buf(w84, k74);
and(x84, o75, e74, k39, j74);
not(y84, m74);
buf(z84, n74);
and(a85, o74, m75, n74);
buf(b85, n74);
and(c85, o74, n74);
and(d85, n74, m75, n39, i74);
and(e85, n74, m75, f74, n39, i74);
and(f85, n74, m75, n39, i74);
and(g85, n74, m75, n39);
and(h85, n74, n39);
and(i85, n74, m75, n39);
and(j85, k74, n75, o39, h74);
and(k85, k74, n75, g74, o39, h74);
and(l85, k74, o39);
and(m85, k74, n75, o39);
buf(n85, o74);
buf(o85, o74);
and(p85, l74, o75, e74, q39, j74);
not(q85, p74);
buf(r85, r74);
not(s85, s74);
not(t85, t74);
buf(u85, u74);
buf(v85, u74);
not(w85, v74);
not(x85, w74);
buf(y85, x74);
buf(z85, x74);
not(t_964, d75);
not(t_965, y74);
or(a86, t_964, t_965);
not(t_966, d77);
not(t_967, z74);
or(b86, t_966, t_967);
not(t_968, b75);
not(t_969, a75);
or(c86, t_968, t_969);
not(t_970, b77);
not(t_971, c75);
or(d86, t_970, t_971);
not(t_972, r75);
not(t_973, e75);
or(e86, t_972, t_973);
not(t_974, y76);
not(t_975, f75);
or(f86, t_974, t_975);
not(t_976, t75);
not(t_977, g75);
or(g86, t_976, t_977);
not(t_978, i77);
not(t_979, h75);
or(h86, t_978, t_979);
not(t_980, a76);
not(t_981, i75);
or(i86, t_980, t_981);
not(t_982, h77);
not(t_983, d65);
or(j86, t_982, t_983);
not(t_984, g76);
not(t_985, j75);
or(k86, t_984, t_985);
not(t_986, g65);
not(t_987, k75);
or(l86, t_986, t_987);
not(t_988, i65);
not(t_989, l75);
or(m86, t_988, t_989);
and(n86, i74, c41);
and(o86, i74, c41);
and(p86, i74, f74, c41);
and(q86, h74, d41);
and(r86, h74, g74, d41);
buf(s86, m75);
buf(t86, m75);
buf(u86, n75);
and(v86, j74, e74, e41);
not(t_990, l76);
not(t_991, p75);
or(w86, t_990, t_991);
not(t_992, r65);
not(t_993, c78);
or(x86, t_992, t_993);
not(t_994, q75);
not(t_995, a78);
or(y86, t_994, t_995);
not(t_996, x76);
not(t_997, s75);
or(z86, t_996, t_997);
not(t_998, x75);
not(t_999, u75);
or(a87, t_998, t_999);
not(t_1000, e76);
not(t_1001, v75);
or(b87, t_1000, t_1001);
not(t_1002, z75);
not(t_1003, w75);
or(c87, t_1002, t_1003);
not(t_1004, t76);
not(t_1005, y75);
or(d87, t_1004, t_1005);
not(t_1006, c76);
not(t_1007, b76);
or(e87, t_1006, t_1007);
not(t_1008, n66);
not(t_1009, g77);
or(f87, t_1008, t_1009);
not(t_1010, q66);
not(t_1011, q77);
or(g87, t_1010, t_1011);
not(t_1012, s76);
not(t_1013, d76);
or(h87, t_1012, t_1013);
not(t_1014, u76);
not(t_1015, f76);
or(i87, t_1014, t_1015);
not(t_1016, w66);
not(t_1017, v76);
or(j87, t_1016, t_1017);
not(t_1018, h76);
not(t_1019, j76);
or(k87, t_1018, t_1019);
not(t_1020, z66);
not(t_1021, z77);
or(l87, t_1020, t_1021);
not(t_1022, b67);
not(t_1023, b78);
or(m87, t_1022, t_1023);
not(t_1024, k76);
not(t_1025, i76);
or(n87, t_1024, t_1025);
not(t_1026, e67);
not(t_1027, w77);
or(o87, t_1026, t_1027);
not(p87, m76);
not(t_1028, n76);
not(t_1029, e77);
or(q87, t_1028, t_1029);
not(r87, o76);
not(t_1030, p67);
not(t_1031, p76);
or(s87, t_1030, t_1031);
not(t_1032, q76);
not(t_1033, r76);
or(t87, t_1032, t_1033);
not(t_1034, s67);
not(t_1035, f77);
or(u87, t_1034, t_1035);
not(t_1036, v67);
not(t_1037, u77);
or(v87, t_1036, t_1037);
not(t_1038, w76);
not(t_1039, z76);
or(w87, t_1038, t_1039);
not(t_1040, a77);
not(t_1041, c77);
or(x87, t_1040, t_1041);
not(y87, j77);
not(t_1042, q68);
not(t_1043, k77);
or(z87, t_1042, t_1043);
not(t_1044, z73);
not(t_1045, a31);
or(a88, t_1044, t_1045);
not(b88, o77);
not(t_1046, y73);
not(t_1047, d25);
or(c88, t_1046, t_1047);
not(d88, r77);
not(t_1048, t77);
not(t_1049, s77);
or(e88, t_1048, t_1049);
not(t_1050, y77);
not(t_1051, v77);
or(f88, t_1050, t_1051);
not(g88, x77);
not(t_1052, d78);
not(t_1053, o69);
or(h88, t_1052, t_1053);
not(i88, e78);
not(t_1054, j78);
not(t_1055, s43);
or(j88, t_1054, t_1055);
not(t_1056, i78);
not(t_1057, t43);
or(k88, t_1056, t_1057);
not(l88, k78);
buf(m88, l78);
buf(n88, l78);
not(o88, m78);
not(p88, o78);
not(q88, p78);
not(r88, q78);
not(s88, r78);
buf(t88, s78);
buf(u88, s78);
not(v88, t78);
not(w88, u78);
and(x88, q59, b84);
and(y88, d79, c79, a79, x78);
buf(z88, x78);
buf(a89, x78);
buf(b89, y78);
buf(c89, y78);
and(d89, z78, e79, b79, y78);
and(e89, y78, b46);
and(f89, x78, c46);
buf(g89, z78);
buf(h89, z78);
and(i89, e79, b79, z78);
buf(j89, a79);
and(k89, d79, c79, a79);
buf(l89, a79);
and(m89, z78, y78, d46);
and(n89, z78, d46);
and(o89, z78, d46);
and(p89, a79, e46);
and(q89, a79, x78, e46);
and(r89, a79, e46);
buf(s89, b79);
buf(t89, b79);
and(u89, e79, b79);
and(v89, d79, c79);
buf(w89, c79);
buf(x89, c79);
and(y89, b79, y78, f46, z78);
and(z89, f46, b79, z78);
and(a90, b79, f46, z78);
and(b90, b79, f46);
and(c90, b79, f46);
and(d90, c79, g46, a79);
and(e90, c79, x78, g46, a79);
and(f90, c79, g46, a79);
and(g90, c79, g46);
buf(h90, d79);
buf(i90, d79);
not(j90, e79);
buf(k90, f79);
buf(l90, f79);
and(m90, o79, l79, j79, i79, f79);
and(n90, h79, n79, k79, g79, m79);
buf(o90, g79);
and(p90, g79, l46);
and(q90, f79, m46);
buf(r90, h79);
buf(s90, i79);
and(t90, o79, j79, i79, l79);
buf(u90, i79);
and(v90, h79, n46);
and(w90, h79, g79, n46);
and(x90, i79, o46);
and(y90, i79, o46);
and(z90, i79, f79, o46);
buf(a91, j79);
buf(b91, j79);
and(c91, o79, j79, l79);
buf(d91, k79);
and(e91, k79, p46, h79);
and(f91, k79, g79, p46, h79);
and(g91, p46, k79);
and(h91, j79, q46, i79);
and(i91, j79, q46, i79);
and(j91, j79, f79, q46, i79);
and(k91, j79, q46);
and(l91, j79, q46);
buf(m91, l79);
buf(n91, l79);
and(o91, o79, l79);
buf(p91, m79);
and(q91, m79, k79, r46, h79);
and(r91, m79, k79, g79, r46, h79);
and(s91, m79, r46);
and(t91, m79, k79, r46);
and(u91, l79, j79, s46, i79);
and(v91, l79, j79, f79, s46, i79);
and(w91, l79, j79, s46, i79);
and(x91, l79, j79, s46);
and(y91, l79, s46);
and(z91, l79, j79, s46);
buf(a92, n79);
buf(b92, o79);
buf(c92, o79);
and(d92, v79, t79, s79, p79);
buf(e92, p79);
buf(f92, p79);
buf(g92, q79);
buf(h92, q79);
and(i92, r79, w79, u79, q79);
and(j92, q79, w46);
and(k92, p79, x46);
buf(l92, r79);
buf(m92, r79);
and(n92, w79, u79, r79);
buf(o92, s79);
and(p92, v79, t79, s79);
buf(q92, s79);
and(r92, r79, q79, y46);
and(s92, r79, y46);
and(t92, r79, y46);
and(u92, s79, z46);
and(v92, s79, p79, z46);
and(w92, s79, z46);
and(x92, v79, t79);
buf(y92, t79);
buf(z92, t79);
buf(a93, u79);
buf(b93, u79);
and(c93, w79, u79);
and(d93, u79, q79, a47, r79);
and(e93, a47, u79, r79);
and(f93, u79, a47, r79);
and(g93, u79, a47);
and(h93, u79, a47);
and(i93, t79, b47, s79);
and(j93, t79, p79, b47, s79);
and(k93, t79, b47, s79);
and(l93, t79, b47);
buf(m93, v79);
buf(n93, v79);
not(o93, w79);
buf(p93, x79);
buf(q93, y79);
buf(r93, y79);
and(s93, x79, g47);
and(t93, y79, h47);
buf(u93, z79);
buf(v93, z79);
buf(w93, a80);
and(x93, a80, i47);
and(y93, a80, x79, i47);
and(z93, z79, j47);
and(a94, z79, j47);
and(b94, z79, y79, j47);
buf(c94, b80);
buf(d94, c80);
buf(e94, c80);
and(f94, b80, k47, a80);
and(g94, b80, x79, k47, a80);
and(h94, k47, b80);
and(i94, c80, l47, z79);
and(j94, c80, l47, z79);
and(k94, c80, y79, l47, z79);
and(l94, c80, l47);
and(m94, c80, l47);
buf(n94, d80);
buf(o94, d80);
buf(p94, e80);
or(q94, w81, c81, n80, t36);
not(t_1058, d81);
not(t_1059, r72);
or(r94, t_1058, t_1059);
and(s94, g80, z81);
and(t94, h80, c82);
not(u94, i80);
not(v94, j80);
or(w94, l81, x80, s80, w36);
or(x94, o81, z80, o80, x36);
not(y94, k80);
not(z94, l80);
and(a95, m80, d82);
not(t_1060, b37);
not(t_1061, b81);
not(t_1062, p81);
and(b95, t_1060, t_1061, t_1062);
or(c95, r80, q81, a81, b37);
not(d95, p80);
not(e95, q80);
not(t_1063, c37);
not(t_1064, w80);
not(t_1065, m81);
and(f95, t_1063, t_1064, t_1065);
or(g95, u80, k81, y80, c37);
not(h95, t80);
not(i95, v80);
or(j95, n81, d37);
not(t_1066, e37);
not(t_1067, s81);
and(k95, t_1066, t_1067);
or(l95, j81, r81, e37);
not(t_1068, f80);
not(t_1069, z72);
or(m95, t_1068, t_1069);
not(n95, f81);
not(o95, g81);
not(p95, h81);
not(q95, i81);
not(t_1070, w61);
not(t_1071, h81);
or(r95, t_1070, t_1071);
not(t_1072, b48);
not(t_1073, i81);
or(s95, t_1072, t_1073);
not(t95, u81);
not(u95, v81);
or(v95, w83, j83, r82, l82, p37);
and(w95, s82, x83, x81);
not(x95, x81);
not(y95, y81);
or(z95, l83, z82, o82, f82, s37);
not(a96, a82);
not(b96, b82);
not(c96, c82);
or(d96, r83, d83, q82, g82, t37);
not(e96, e82);
not(t_1074, u37);
not(t_1075, m82);
not(t_1076, x82);
not(t_1077, m83);
and(f96, t_1074, t_1075, t_1076, t_1077);
or(g96, j82, k83, y82, n82, u37);
not(h96, h82);
not(i96, i82);
not(j96, k82);
not(t_1078, z37);
not(t_1079, a83);
not(t_1080, p83);
and(k96, t_1078, t_1079, t_1080);
or(l96, v82, n83, b83, z37);
and(m96, m73, u73, y81);
not(n96, t82);
not(o96, u82);
not(p96, w82);
or(q96, o83, e38);
not(r96, f83);
not(s96, g83);
not(t96, h83);
not(u96, u83);
not(v96, v83);
not(w96, y83);
and(x96, k49, f84);
and(y96, n49, e84);
or(z96, e85, q84, p86, h84, y38);
or(a97, k85, u84, r86, i84, z38);
or(b97, p85, x84, v86, n84, a39);
and(c97, y84, q85, z83);
not(d97, z83);
not(e97, a84);
not(f97, c84);
not(g97, d84);
not(h97, e84);
not(i97, g84);
not(t_1081, d39);
not(t_1082, n86);
not(t_1083, o84);
not(t_1084, f85);
and(j97, t_1081, t_1082, t_1083, t_1084);
or(k97, l84, d85, p84, o86, d39);
not(l97, j84);
not(m97, k84);
not(n97, m84);
or(o97, h85, i39);
not(p97, w84);
and(q97, m74, p74, a84);
not(r97, z84);
not(s97, b85);
not(t97, n85);
not(u97, o85);
not(v97, r85);
and(w97, t74, s74, u85);
and(x97, t85, s85, v85);
not(y97, u85);
not(z97, v85);
and(a98, w74, v74, y85);
and(b98, x85, w85, z85);
not(c98, y85);
not(d98, z85);
not(e98, a86);
and(f98, d86, z86, k51, f86);
and(g98, b86, d86, f86, z86);
not(h98, c86);
and(i98, f86, z86, s51);
not(j98, e86);
and(k98, z86, y51);
not(l98, g86);
buf(m98, h86);
buf(n98, h86);
and(o98, f87, e52);
and(p98, k86, b87, d87, i86, f87);
buf(q98, j86);
buf(r98, j86);
and(s98, b87, d87, f87, h52, i86);
not(t98, l86);
not(u98, m86);
not(t_1085, c41);
not(t_1086, r84);
not(t_1087, i85);
and(v98, t_1085, t_1086, t_1087);
or(w98, a85, g85, s84, c41);
not(x98, s86);
not(y98, t86);
not(z98, u86);
and(a99, h88, o87, l87, m87, w86);
buf(b99, x86);
buf(c99, x86);
buf(d99, y86);
buf(e99, y86);
not(f99, a87);
and(g99, d87, f87, i53, i86);
not(h99, c87);
and(i99, i86, f87, p53);
buf(j99, e87);
buf(k99, e87);
and(l99, g87, v87, u87, s87);
not(m99, h87);
not(n99, i87);
not(o99, j87);
not(p99, k87);
buf(q99, n87);
buf(r99, n87);
not(s99, q87);
not(t_1088, d88);
not(t_1089, o76);
or(t99, t_1088, t_1089);
not(u99, t87);
not(v99, w87);
not(w99, x87);
and(x99, s87, l55);
not(y99, z87);
not(t_1090, a88);
not(t_1091, m77);
or(z99, t_1090, t_1091);
not(t_1092, c88);
not(t_1093, p77);
or(a100, t_1092, t_1093);
and(b100, v87, s87, c56, u87);
not(t_1094, r87);
not(t_1095, r77);
or(c100, t_1094, t_1095);
not(d100, e88);
and(e100, u87, s87, l56);
not(f100, f88);
and(g100, l87, w86, r56, m87);
and(h100, m87, w86, y56);
and(i100, w86, d57);
and(j100, o87, l87, w86, g57, m87);
and(k100, e80, b80, p69, a80);
and(l100, e80, b80, x79, p69, a80);
and(m100, e80, p69);
and(n100, e80, b80, p69);
and(o100, d80, c80, q69, z79);
and(p100, d80, c80, y79, q69, z79);
and(q100, d80, c80, q69, z79);
and(r100, d80, c80, q69);
and(s100, d80, q69);
and(t100, d80, c80, q69);
not(t_1096, j88);
not(t_1097, f78);
or(u100, t_1096, t_1097);
not(t_1098, k88);
not(t_1099, h78);
or(v100, t_1098, t_1099);
and(w100, m78, k78, n88);
and(x100, o88, l88, m88);
not(y100, m88);
not(z100, n88);
not(t_1100, q88);
not(t_1101, o78);
or(a101, t_1100, t_1101);
not(t_1102, p88);
not(t_1103, p78);
or(b101, t_1102, t_1103);
not(t_1104, s88);
not(t_1105, q78);
or(c101, t_1104, t_1105);
not(t_1106, r88);
not(t_1107, r78);
or(d101, t_1106, t_1107);
and(e101, v88, w88, t88);
not(f101, t88);
not(g101, u88);
and(h101, t78, u78, u88);
and(i101, q59, b97);
and(j101, x6, u100);
and(k101, x6, u100, e80);
and(l101, x6, u100, b80, e80);
and(m101, x6, u100, b80, e80, a80);
or(n101, y89, m89, e89, z45);
or(o101, e90, q89, f89, a46);
and(p101, y88, m90);
not(q101, z88);
not(r101, a89);
not(s101, b89);
not(t101, c89);
and(u101, d89, n90);
not(t_1108, b46);
not(t_1109, o89);
not(t_1110, z89);
and(v101, t_1108, t_1109, t_1110);
or(w101, i89, a90, n89, b46);
not(t_1111, c46);
not(t_1112, p89);
not(t_1113, f90);
and(x101, t_1111, t_1112, t_1113);
or(y101, k89, d90, r89, c46);
not(z101, g89);
not(a102, h89);
not(b102, j89);
not(c102, l89);
not(t_1114, d46);
not(t_1115, c90);
and(d102, t_1114, t_1115);
or(e102, u89, b90, d46);
or(f102, g90, e46);
not(g102, s89);
not(h102, t89);
not(i102, w89);
not(j102, x89);
not(t_1116, k71);
not(t_1117, s89);
or(k102, t_1116, t_1117);
not(l102, h90);
not(m102, i90);
not(t_1118, c60);
not(t_1119, t89);
or(n102, t_1118, t_1119);
or(o102, r91, f91, w90, p90, j46);
or(p102, v91, j91, z90, q90, k46);
not(q102, k90);
not(r102, l90);
not(s102, m90);
not(t102, o90);
not(t_1120, m46);
not(t_1121, x90);
not(t_1122, h91);
not(t_1123, w91);
and(u102, t_1120, t_1121, t_1122, t_1123);
or(v102, t90, u91, i91, y90, m46);
not(w102, r90);
not(x102, s90);
not(y102, u90);
not(t_1124, o46);
not(t_1125, k91);
not(t_1126, z91);
and(z102, t_1124, t_1125, t_1126);
or(a103, c91, x91, l91, o46);
not(b103, a91);
not(c103, b91);
not(d103, d91);
or(e103, y91, q46);
not(f103, m91);
not(g103, n91);
not(h103, p91);
not(i103, a92);
not(j103, b92);
not(k103, c92);
or(l103, d93, r92, j92, u46);
or(m103, j93, v92, k92, v46);
not(n103, d92);
not(o103, e92);
not(p103, f92);
not(q103, g92);
not(r103, h92);
not(s103, i92);
not(t_1127, w46);
not(t_1128, t92);
not(t_1129, e93);
and(t103, t_1127, t_1128, t_1129);
or(u103, n92, f93, s92, w46);
not(t_1130, x46);
not(t_1131, u92);
not(t_1132, k93);
and(v103, t_1130, t_1131, t_1132);
or(w103, p92, i93, w92, x46);
not(x103, l92);
not(y103, m92);
not(z103, o92);
not(a104, q92);
not(t_1133, y46);
not(t_1134, h93);
and(b104, t_1133, t_1134);
or(c104, c93, g93, y46);
or(d104, l93, z46);
not(e104, y92);
not(f104, z92);
not(g104, a93);
not(h104, b93);
not(t_1135, f72);
not(t_1136, a93);
or(i104, t_1135, t_1136);
not(j104, m93);
not(k104, n93);
not(t_1137, a61);
not(t_1138, b93);
or(l104, t_1137, t_1138);
or(m104, l100, g94, y93, s93, e47);
or(n104, p100, k94, b94, t93, f47);
and(o104, a80, u100, b80, x79, e80);
not(p104, p93);
not(q104, q93);
not(r104, r93);
and(s104, v100, d80, c80, z79, y79);
not(t_1139, h47);
not(t_1140, z93);
not(t_1141, i94);
not(t_1142, q100);
and(t104, t_1139, t_1140, t_1141, t_1142);
not(u104, u93);
and(v104, v100, c80, z79, d80);
not(w104, v93);
not(x104, w93);
not(t_1143, j47);
not(t_1144, l94);
not(t_1145, t100);
and(y104, t_1143, t_1144, t_1145);
not(z104, c94);
not(a105, d94);
not(b105, e94);
and(c105, v100, c80, d80);
or(d105, s100, l47);
not(e105, n94);
not(f105, o94);
and(g105, v100, d80);
not(h105, p94);
not(t_1146, r94);
not(t_1147, m95);
or(i105, t_1146, t_1147);
and(j105, g80, v95);
and(k105, h80, z95);
not(t_1148, y94);
not(t_1149, c95);
or(l105, t_1148, t_1149);
not(t_1150, z94);
not(t_1151, b95);
or(m105, t_1150, t_1151);
and(n105, d96, m80);
not(o105, b95);
not(p105, c95);
not(t_1152, d95);
not(t_1153, k95);
or(q105, t_1152, t_1153);
not(t_1154, e95);
not(t_1155, l95);
or(r105, t_1154, t_1155);
not(s105, f95);
not(t105, g95);
not(u105, j95);
not(v105, k95);
not(w105, l95);
or(x105, e81, j95);
not(t_1156, p95);
not(t_1157, z47);
or(y105, t_1156, t_1157);
not(t_1158, q95);
not(t_1159, k37);
or(z105, t_1158, t_1159);
not(a106, z95);
not(b106, f96);
not(c106, g96);
not(d106, k96);
not(e106, l96);
and(f106, x83, m73, y95);
not(g106, q96);
or(h106, i83, q96);
not(t_1160, r62);
not(t_1161, k96);
or(i106, t_1160, t_1161);
not(t_1162, x48);
not(t_1163, l96);
or(j106, t_1162, t_1163);
and(k106, u73, s82, x95);
not(t_1164, z62);
not(t_1165, z99);
or(l106, t_1164, t_1165);
not(t_1166, b74);
not(t_1167, a100);
or(m106, t_1166, t_1167);
and(n106, a97, k49);
and(o106, n49, z96);
not(p106, z96);
not(q106, b97);
not(r106, j97);
not(s106, k97);
not(t106, o97);
and(u106, q85, m74, e97);
or(v106, c85, o97);
not(t_1168, t63);
not(t_1169, v98);
or(w106, t_1168, t_1169);
not(t_1170, h50);
not(t_1171, w98);
or(x106, t_1170, t_1171);
and(y106, p74, y84, d97);
and(z106, s74, t85, z97);
and(a107, s85, t74, y97);
and(b107, v74, x85, d98);
and(c107, w85, w74, c98);
not(t_1172, l98);
not(t_1173, a86);
or(d107, t_1172, t_1173);
and(e107, g98, a99);
not(f107, g98);
not(t_1174, j98);
not(t_1175, c86);
or(g107, t_1174, t_1175);
not(t_1176, h98);
not(t_1177, e86);
or(h107, t_1176, t_1177);
not(t_1178, e98);
not(t_1179, g86);
or(i107, t_1178, t_1179);
and(j107, f99, u98, m98);
not(k107, m98);
not(l107, n98);
and(m107, l99, p98);
and(n107, h99, t98, q98);
not(o107, q98);
not(p107, r98);
and(q107, c87, l86, r98);
and(r107, a87, m86, n98);
not(s107, v98);
not(t107, w98);
or(u107, j100, g100, h100, i100, u52);
not(v107, b99);
not(w107, c99);
not(x107, d99);
and(y107, f100, y99, e99);
not(z107, e99);
or(a108, f98, i98, k98, d53);
not(t_1180, w0);
not(t_1181, a99);
or(b108, t_1180, t_1181);
not(c108, j99);
and(d108, n99, o99, k99);
not(e108, k99);
not(f108, l99);
not(t_1182, u99);
not(t_1183, h87);
or(g108, t_1182, t_1183);
and(h108, i87, j87, j99);
not(i108, q99);
not(j108, r99);
and(k108, k87, m76, r99);
and(l108, p99, p87, q99);
not(t_1184, d100);
not(t_1185, q87);
or(m108, t_1184, t_1185);
or(n108, b100, e100, x99, o54);
not(t_1186, t99);
not(t_1187, c100);
or(o108, t_1186, t_1187);
not(t_1188, m99);
not(t_1189, t87);
or(p108, t_1188, t_1189);
not(t_1190, w99);
not(t_1191, w87);
or(q108, t_1190, t_1191);
not(t_1192, v99);
not(t_1193, x87);
or(r108, t_1192, t_1193);
or(s108, s98, g99, i99, o98, o55);
and(t108, x77, j77, c99);
and(u108, g88, y87, b99);
and(v108, f88, z87, d99);
not(w108, z99);
not(x108, a100);
not(t_1194, s99);
not(t_1195, e88);
or(y108, t_1194, t_1195);
buf(z108, u100);
buf(a109, v100);
buf(b109, v100);
and(c109, k78, o88, y100);
and(d109, l88, m78, z100);
not(t_1196, a101);
not(t_1197, b101);
or(e109, t_1196, t_1197);
not(t_1198, d101);
not(t_1199, c101);
or(f109, t_1198, t_1199);
and(g109, w88, t78, g101);
and(h109, u78, v88, f101);
not(t_1200, d16);
not(t_1201, z108);
or(i109, t_1200, t_1201);
not(t_1202, x6);
not(t_1203, s104);
or(j109, t_1202, t_1203);
and(k109, o104, x6);
and(l109, y88, p102);
not(t_1204, s101);
not(t_1205, w101);
or(m109, t_1204, t_1205);
not(t_1206, t101);
not(t_1207, v101);
or(n109, t_1206, t_1207);
and(o109, o102, d89);
not(p109, v101);
not(q109, w101);
not(r109, x101);
not(s109, y101);
not(t_1208, z101);
not(t_1209, d102);
or(t109, t_1208, t_1209);
not(t_1210, a102);
not(t_1211, e102);
or(u109, t_1210, t_1211);
not(v109, d102);
not(w109, e102);
not(x109, f102);
or(y109, v89, f102);
not(t_1212, g102);
not(t_1213, x59);
or(z109, t_1212, t_1213);
not(t_1214, h102);
not(t_1215, i46);
or(a110, t_1214, t_1215);
not(b110, p102);
not(c110, u102);
not(d110, v102);
not(e110, z102);
not(f110, a103);
not(g110, e103);
or(h110, o91, e103);
not(t_1216, w71);
not(t_1217, z102);
or(i110, t_1216, t_1217);
not(t_1218, n60);
not(t_1219, a103);
or(j110, t_1218, t_1219);
not(k110, l103);
not(l110, m103);
and(m110, d92, n104);
and(n110, d92, s104);
not(t_1220, q103);
not(t_1221, u103);
or(o110, t_1220, t_1221);
not(t_1222, r103);
not(t_1223, t103);
or(p110, t_1222, t_1223);
and(q110, i92, o104);
and(r110, m104, i92);
not(s110, t103);
not(t110, u103);
not(u110, v103);
not(v110, w103);
not(t_1224, x103);
not(t_1225, b104);
or(w110, t_1224, t_1225);
not(t_1226, y103);
not(t_1227, c104);
or(x110, t_1226, t_1227);
not(y110, b104);
not(z110, c104);
not(a111, d104);
or(b111, x92, d104);
not(t_1228, g104);
not(t_1229, v60);
or(c111, t_1228, t_1229);
not(t_1230, h104);
not(t_1231, d47);
or(d111, t_1230, t_1231);
not(e111, n104);
not(f111, s104);
or(g111, m101, k100, f94, x93, g47);
not(h111, t104);
or(i111, v104, o100, j94, a94, h47);
or(j111, l101, n100, h94, i47);
not(k111, y104);
or(l111, c105, r100, m94, j47);
or(m111, k101, m100, k47);
or(n111, g105, d105);
not(o111, d105);
or(p111, j105, q94);
not(q111, i105);
or(r111, k105, w94);
or(s111, n105, x94);
not(t_1232, p105);
not(t_1233, k80);
or(t111, t_1232, t_1233);
not(t_1234, o105);
not(t_1235, l80);
or(u111, t_1234, t_1235);
not(t_1236, v105);
not(t_1237, p80);
or(v111, t_1236, t_1237);
not(t_1238, w105);
not(t_1239, q80);
or(w111, t_1238, t_1239);
not(x111, u105);
not(y111, x105);
not(t_1240, v61);
not(t_1241, u105);
or(z111, t_1240, t_1241);
not(t_1242, y105);
not(t_1243, r95);
or(a112, t_1242, t_1243);
not(t_1244, z105);
not(t_1245, s95);
or(b112, t_1244, t_1245);
not(t_1246, c48);
not(t_1247, x105);
or(c112, t_1246, t_1247);
not(t_1248, k106);
not(t_1249, w95);
and(d112, t_1248, t_1249);
and(e112, a106, c96);
not(t_1250, f106);
not(t_1251, m96);
and(f112, t_1250, t_1251);
not(g112, g106);
not(h112, h106);
not(t_1252, d106);
not(t_1253, w48);
or(i112, t_1252, t_1253);
not(t_1254, e106);
not(t_1255, l38);
or(j112, t_1254, t_1255);
not(t_1256, w108);
not(t_1257, f49);
or(k112, t_1256, t_1257);
or(l112, o106, g49);
not(t_1258, x108);
not(t_1259, b63);
or(m112, t_1258, t_1259);
or(n112, n106, h49);
not(t_1260, y106);
not(t_1261, c97);
and(o112, t_1260, t_1261);
and(p112, p106, h97);
not(q112, t106);
not(t_1262, u106);
not(t_1263, q97);
and(r112, t_1262, t_1263);
not(s112, v106);
not(t_1264, s107);
not(t_1265, g50);
or(t112, t_1264, t_1265);
not(t_1266, t107);
not(t_1267, p39);
or(u112, t_1266, t_1267);
not(t_1268, a107);
not(t_1269, w97);
and(v112, t_1268, t_1269);
not(t_1270, z106);
not(t_1271, x97);
and(w112, t_1270, t_1271);
not(t_1272, c107);
not(t_1273, a98);
and(x112, t_1272, t_1273);
not(t_1274, b107);
not(t_1275, b98);
and(y112, t_1274, t_1275);
not(t_1276, i107);
not(t_1277, d107);
or(z112, t_1276, t_1277);
and(a113, g98, u107);
not(t_1278, h107);
not(t_1279, g107);
or(b113, t_1278, t_1279);
and(c113, l86, h99, o107);
and(d113, m86, f99, k107);
not(e113, u107);
not(f113, a108);
and(g113, u98, a87, l107);
and(h113, t98, c87, p107);
and(i113, w0, e107, m107, s94, x88);
and(j113, w0, e107, m107, s94);
and(k113, w0, e107, m107, s94, x88);
and(l113, l99, s108);
not(t_1280, p108);
not(t_1281, g108);
or(m113, t_1280, t_1281);
and(n113, o99, i87, c108);
and(o113, j87, n99, e108);
and(p113, p87, k87, j108);
and(q113, m76, p99, i108);
not(t_1282, m108);
not(t_1283, y108);
or(r113, t_1282, t_1283);
not(s113, n108);
not(t113, o108);
not(t_1284, q108);
not(t_1285, r108);
or(u113, t_1284, t_1285);
not(v113, s108);
and(w113, j77, g88, v107);
and(x113, z87, f100, z107);
or(y113, i101, s68);
and(z113, y99, f88, x107);
and(a114, y87, x77, w107);
or(b114, j101, p69);
not(t_1286, i88);
not(t_1287, y104);
or(c114, t_1286, t_1287);
not(d114, z108);
not(e114, a109);
not(f114, b109);
not(t_1288, d109);
not(t_1289, w100);
and(g114, t_1288, t_1289);
not(t_1290, c109);
not(t_1291, x100);
and(h114, t_1290, t_1291);
not(i114, e109);
not(j114, f109);
not(t_1292, h109);
not(t_1293, e101);
and(k114, t_1292, t_1293);
not(t_1294, g109);
not(t_1295, h101);
and(l114, t_1294, t_1295);
and(m114, p111, x88);
and(n114, p111, x88);
not(t_1296, d114);
not(t_1297, m13);
or(o114, t_1296, t_1297);
and(p114, x6, q110, u101);
and(q114, x6, q110, u101, a95);
and(r114, e111, j109);
and(s114, x6, n110, p101);
and(t114, x6, n110, p101, t94);
and(u114, x6, n110, p101, t94, y96);
and(v114, x6, q110, u101, a95, x96);
or(w114, o109, n101);
or(x114, l109, o101);
not(t_1298, q109);
not(t_1299, b89);
or(y114, t_1298, t_1299);
not(t_1300, p109);
not(t_1301, c89);
or(z114, t_1300, t_1301);
not(t_1302, v109);
not(t_1303, g89);
or(a115, t_1302, t_1303);
not(t_1304, w109);
not(t_1305, h89);
or(b115, t_1304, t_1305);
not(c115, x109);
not(d115, y109);
not(t_1306, z109);
not(t_1307, k102);
or(e115, t_1306, t_1307);
not(t_1308, l71);
not(t_1309, x109);
or(f115, t_1308, t_1309);
not(t_1310, z59);
not(t_1311, y109);
or(g115, t_1310, t_1311);
not(t_1312, a110);
not(t_1313, n102);
or(h115, t_1312, t_1313);
and(i115, b110, s102);
not(j115, g110);
not(k115, h110);
not(t_1314, e110);
not(t_1315, l60);
or(l115, t_1314, t_1315);
not(t_1316, f110);
not(t_1317, t46);
or(m115, t_1316, t_1317);
or(n115, r110, l103);
or(o115, m110, m103);
not(t_1318, n103);
not(t_1319, l110);
or(p115, t_1318, t_1319);
not(t_1320, t110);
not(t_1321, g92);
or(q115, t_1320, t_1321);
not(t_1322, s110);
not(t_1323, h92);
or(r115, t_1322, t_1323);
not(t_1324, s103);
not(t_1325, k110);
or(s115, t_1324, t_1325);
not(t_1326, y110);
not(t_1327, l92);
or(t115, t_1326, t_1327);
not(t_1328, z110);
not(t_1329, m92);
or(u115, t_1328, t_1329);
not(v115, a111);
not(w115, b111);
not(t_1330, c111);
not(t_1331, i104);
or(x115, t_1330, t_1331);
not(t_1332, g72);
not(t_1333, a111);
or(y115, t_1332, t_1333);
not(t_1334, x60);
not(t_1335, b111);
or(z115, t_1334, t_1335);
not(t_1336, d111);
not(t_1337, l104);
or(a116, t_1336, t_1337);
or(b116, k109, m104);
and(c116, e111, f111);
not(t_1338, p104);
not(t_1339, g111);
or(d116, t_1338, t_1339);
not(e116, g111);
not(f116, i111);
not(t_1340, x104);
not(t_1341, j111);
or(g116, t_1340, t_1341);
not(h116, j111);
not(i116, l111);
not(t_1342, z104);
not(t_1343, m111);
or(j116, t_1342, t_1343);
not(k116, m111);
not(l116, n111);
not(m116, o111);
not(t_1344, h105);
not(t_1345, b114);
or(n116, t_1344, t_1345);
not(t_1346, l105);
not(t_1347, t111);
or(o116, t_1346, t_1347);
not(t_1348, m105);
not(t_1349, u111);
or(p116, t_1348, t_1349);
not(t_1350, q105);
not(t_1351, v111);
or(q116, t_1350, t_1351);
not(t_1352, r105);
not(t_1353, w111);
or(r116, t_1352, t_1353);
not(t_1354, x111);
not(t_1355, y47);
or(s116, t_1354, t_1355);
not(t116, b112);
not(t_1356, y111);
not(t_1357, l37);
or(u116, t_1356, t_1357);
not(t_1358, f112);
not(t_1359, d112);
or(v116, t_1358, t_1359);
not(w116, e112);
not(t_1360, i112);
not(t_1361, i106);
or(x116, t_1360, t_1361);
not(t_1362, j112);
not(t_1363, j106);
or(y116, t_1362, t_1363);
not(t_1364, l106);
not(t_1365, k112);
or(z116, t_1364, t_1365);
not(t_1366, m106);
not(t_1367, m112);
or(a117, t_1366, t_1367);
and(b117, s111, x96);
and(c117, r111, y96);
not(t_1368, r112);
not(t_1369, o112);
or(d117, t_1368, t_1369);
not(e117, p112);
not(t_1370, t112);
not(t_1371, w106);
or(f117, t_1370, t_1371);
not(t_1372, u112);
not(t_1373, x106);
or(g117, t_1372, t_1373);
not(t_1374, v112);
not(t_1375, w112);
or(h117, t_1374, t_1375);
not(t_1376, x112);
not(t_1377, y112);
or(i117, t_1376, t_1377);
not(j117, z112);
not(t_1378, f107);
not(t_1379, f113);
or(k117, t_1378, t_1379);
not(l117, b113);
not(t_1380, d113);
not(t_1381, j107);
and(m117, t_1380, t_1381);
not(t_1382, c113);
not(t_1383, n107);
and(n117, t_1382, t_1383);
not(t_1384, h113);
not(t_1385, q107);
and(o117, t_1384, t_1385);
not(t_1386, g113);
not(t_1387, r107);
and(p117, t_1386, t_1387);
not(t_1388, x113);
not(t_1389, y107);
and(q117, t_1388, t_1389);
or(r117, a113, a108);
and(s117, e113, b108);
not(t_1390, o113);
not(t_1391, d108);
and(t117, t_1390, t_1391);
not(t_1392, f108);
not(t_1393, s113);
or(u117, t_1392, t_1393);
not(v117, m113);
not(t_1394, n113);
not(t_1395, h108);
and(w117, t_1394, t_1395);
not(t_1396, p113);
not(t_1397, k108);
and(x117, t_1396, t_1397);
not(t_1398, q113);
not(t_1399, l108);
and(y117, t_1398, t_1399);
not(z117, r113);
or(a118, l113, n108);
not(b118, u113);
not(t_1400, a114);
not(t_1401, t108);
and(c118, t_1400, t_1401);
not(t_1402, w113);
not(t_1403, u108);
and(d118, t_1402, t_1403);
not(t_1404, z113);
not(t_1405, v108);
and(e118, t_1404, t_1405);
not(f118, b114);
not(t_1406, k111);
not(t_1407, e78);
or(g118, t_1406, t_1407);
not(t_1408, g78);
not(t_1409, l111);
or(h118, t_1408, t_1409);
not(t_1410, g114);
not(t_1411, h114);
or(i118, t_1410, t_1411);
not(t_1412, l114);
not(t_1413, k114);
or(j118, t_1412, t_1413);
and(k118, a118, s94, x88);
and(l118, r117, m107, s94, x88);
and(m118, a118, s94, x88);
and(n118, r117, m107, s94, x88);
not(o118, r114);
and(p118, o115, p101);
not(t_1414, m109);
not(t_1415, y114);
or(q118, t_1414, t_1415);
not(t_1416, n109);
not(t_1417, z114);
or(r118, t_1416, t_1417);
and(s118, n115, u101);
not(t_1418, t109);
not(t_1419, a115);
or(t118, t_1418, t_1419);
not(t_1420, u109);
not(t_1421, b115);
or(u118, t_1420, t_1421);
not(t_1422, c115);
not(t_1423, y59);
or(v118, t_1422, t_1423);
not(t_1424, d115);
not(t_1425, h46);
or(w118, t_1424, t_1425);
not(x118, h115);
not(y118, i115);
not(t_1426, l115);
not(t_1427, i110);
or(z118, t_1426, t_1427);
not(t_1428, m115);
not(t_1429, j110);
or(a119, t_1428, t_1429);
and(b119, r114, m103);
not(t_1430, o110);
not(t_1431, q115);
or(c119, t_1430, t_1431);
not(t_1432, p110);
not(t_1433, r115);
or(d119, t_1432, t_1433);
and(e119, s115, b116);
not(t_1434, w110);
not(t_1435, t115);
or(f119, t_1434, t_1435);
not(t_1436, x110);
not(t_1437, u115);
or(g119, t_1436, t_1437);
not(t_1438, v115);
not(t_1439, w60);
or(h119, t_1438, t_1439);
not(t_1440, w115);
not(t_1441, c47);
or(i119, t_1440, t_1441);
and(j119, b116, o93);
not(k119, a116);
not(l119, b116);
not(m119, c116);
not(t_1442, e116);
not(t_1443, p93);
or(n119, t_1442, t_1443);
not(t_1444, h116);
not(t_1445, w93);
or(o119, t_1444, t_1445);
not(t_1446, k116);
not(t_1447, c94);
or(p119, t_1446, t_1447);
not(t_1448, f118);
not(t_1449, p94);
or(q119, t_1448, t_1449);
not(t_1450, q111);
not(t_1451, v116);
or(r119, t_1450, t_1451);
and(s119, a118, s94);
and(t119, r117, m107, s94);
and(u119, x114, t94, y96);
and(v119, o115, p101, t94, y96);
and(w119, x114, t94);
and(x119, o115, p101, t94);
not(y119, p116);
and(z119, w114, a95, x96);
and(a120, n115, u101, a95, x96);
and(b120, w114, a95);
and(c120, n115, u101, a95);
not(d120, q116);
not(t_1452, s116);
not(t_1453, z111);
or(e120, t_1452, t_1453);
not(t_1454, u116);
not(t_1455, c112);
or(f120, t_1454, t_1455);
not(g120, v116);
not(t_1456, g112);
not(t_1457, x116);
or(h120, t_1456, t_1457);
not(t_1458, h112);
not(t_1459, y116);
or(i120, t_1458, t_1459);
not(j120, x116);
not(k120, y116);
not(t_1460, x73);
not(t_1461, d117);
or(l120, t_1460, t_1461);
not(m120, z116);
not(n120, a117);
not(t_1462, f63);
not(t_1463, z116);
or(o120, t_1462, t_1463);
not(t_1464, g63);
not(t_1465, a117);
or(p120, t_1464, t_1465);
not(q120, d117);
not(t_1466, q112);
not(t_1467, f117);
or(r120, t_1466, t_1467);
not(t_1468, s112);
not(t_1469, g117);
or(s120, t_1468, t_1469);
not(t120, f117);
not(u120, g117);
not(v120, h117);
not(w120, i117);
not(t_1470, p117);
not(t_1471, m117);
or(x120, t_1470, t_1471);
not(t_1472, o117);
not(t_1473, n117);
or(y120, t_1472, t_1473);
not(t_1474, e118);
not(t_1475, q117);
or(z120, t_1474, t_1475);
and(a121, s117, a108);
not(b121, s117);
not(t_1476, w117);
not(t_1477, t117);
or(c121, t_1476, t_1477);
not(t_1478, x117);
not(t_1479, y117);
or(d121, t_1478, t_1479);
not(t_1480, c118);
not(t_1481, d118);
or(e121, t_1480, t_1481);
not(t_1482, g118);
not(t_1483, c114);
or(f121, t_1482, t_1483);
not(t_1484, i116);
not(t_1485, r69);
or(g121, t_1484, t_1485);
not(h121, i118);
not(t_1486, n78);
not(t_1487, i118);
or(i121, t_1486, t_1487);
not(t_1488, i114);
not(t_1489, h117);
or(j121, t_1488, t_1489);
not(t_1490, j114);
not(t_1491, i117);
or(k121, t_1490, t_1491);
not(l121, j118);
not(t_1492, v78);
not(t_1493, j118);
or(m121, t_1492, t_1493);
or(n121, p114, s118, w114);
or(o121, s114, p118, x114);
not(p121, r118);
not(q121, t118);
not(t_1494, v118);
not(t_1495, f115);
or(r121, t_1494, t_1495);
not(t_1496, w118);
not(t_1497, g115);
or(s121, t_1496, t_1497);
not(t_1498, j115);
not(t_1499, z118);
or(t121, t_1498, t_1499);
not(t_1500, k115);
not(t_1501, a119);
or(u121, t_1500, t_1501);
not(v121, z118);
not(w121, a119);
and(x121, l103, l119);
and(y121, p115, o118);
not(z121, d119);
not(a122, f119);
and(b122, x115, l119);
not(t_1502, h119);
not(t_1503, y115);
or(c122, t_1502, t_1503);
not(t_1504, i119);
not(t_1505, z115);
or(d122, t_1504, t_1505);
and(e122, w79, l119);
and(f122, b116, c119);
and(g122, b116, g119);
and(h122, b116, k119);
not(t_1506, m116);
not(t_1507, f121);
or(i122, t_1506, t_1507);
or(j122, j113, t119, s119, p111);
not(t_1508, g120);
not(t_1509, i105);
or(k122, t_1508, t_1509);
or(l122, t114, x119, w119, r111);
or(m122, q114, c120, b120, s111);
not(t_1510, s105);
not(t_1511, e120);
or(n122, t_1510, t_1511);
not(t_1512, t105);
not(t_1513, f120);
or(o122, t_1512, t_1513);
not(p122, e120);
not(q122, f120);
not(t_1514, j120);
not(t_1515, g106);
or(r122, t_1514, t_1515);
not(t_1516, k120);
not(t_1517, h106);
or(s122, t_1516, t_1517);
not(t_1518, q120);
not(t_1519, w62);
or(t122, t_1518, t_1519);
not(t_1520, m120);
not(t_1521, r49);
or(u122, t_1520, t_1521);
not(t_1522, n120);
not(t_1523, s49);
or(v122, t_1522, t_1523);
not(t_1524, t120);
not(t_1525, t106);
or(w122, t_1524, t_1525);
not(t_1526, u120);
not(t_1527, v106);
or(x122, t_1526, t_1527);
not(t_1528, j117);
not(t_1529, e121);
or(y122, t_1528, t_1529);
and(z122, k117, b121);
not(t_1530, l117);
not(t_1531, z120);
or(a123, t_1530, t_1531);
not(b123, x120);
not(c123, y120);
not(d123, z120);
not(e123, c121);
not(t_1532, v117);
not(t_1533, c121);
or(f123, t_1532, t_1533);
not(g123, d121);
not(t_1534, z117);
not(t_1535, x120);
or(h123, t_1534, t_1535);
not(t_1536, t113);
not(t_1537, y120);
or(i123, t_1536, t_1537);
not(t_1538, b118);
not(t_1539, d121);
or(j123, t_1538, t_1539);
not(k123, e121);
not(l123, f121);
not(t_1540, g121);
not(t_1541, h118);
or(m123, t_1540, t_1541);
not(t_1542, h121);
not(t_1543, e70);
or(n123, t_1542, t_1543);
not(t_1544, v120);
not(t_1545, e109);
or(o123, t_1544, t_1545);
not(t_1546, w120);
not(t_1547, f109);
or(p123, t_1546, t_1547);
not(t_1548, l121);
not(t_1549, b71);
or(q123, t_1548, t_1549);
buf(r123, n121);
not(s123, o121);
not(t_1550, r109);
not(t_1551, r121);
or(t123, t_1550, t_1551);
not(t_1552, s109);
not(t_1553, s121);
or(u123, t_1552, t_1553);
not(v123, r121);
not(w123, s121);
not(t_1554, v121);
not(t_1555, g110);
or(x123, t_1554, t_1555);
not(t_1556, w121);
not(t_1557, h110);
or(y123, t_1556, t_1557);
or(z123, b119, y121);
or(a124, e119, x121);
not(t_1558, u110);
not(t_1559, c122);
or(b124, t_1558, t_1559);
not(t_1560, v110);
not(t_1561, d122);
or(c124, t_1560, t_1561);
not(d124, c122);
not(e124, d122);
and(f124, z121, l119);
and(g124, a122, l119);
not(t_1562, l116);
not(t_1563, m123);
or(h124, t_1562, t_1563);
not(t_1564, l123);
not(t_1565, o111);
or(i124, t_1564, t_1565);
not(t_1566, r119);
not(t_1567, k122);
or(j124, t_1566, t_1567);
buf(k124, l122);
buf(l124, m122);
not(t_1568, p122);
not(t_1569, f95);
or(m124, t_1568, t_1569);
not(t_1570, q122);
not(t_1571, g95);
or(n124, t_1570, t_1571);
and(o124, d82, n121);
and(p124, n121, w73, p73, q73, j73);
and(q124, n121, w73, p73, q73);
not(t_1572, h120);
not(t_1573, r122);
or(r124, t_1572, t_1573);
and(s124, n121, w73, q73);
not(t_1574, i120);
not(t_1575, s122);
or(t124, t_1574, t_1575);
and(u124, n121, w73);
not(t_1576, l120);
not(t_1577, t122);
or(v124, t_1576, t_1577);
not(t_1578, o120);
not(t_1579, u122);
or(w124, t_1578, t_1579);
not(t_1580, p120);
not(t_1581, v122);
or(x124, t_1580, t_1581);
not(t_1582, j122);
not(t_1583, b84);
or(y124, t_1582, t_1583);
not(t_1584, l122);
not(t_1585, e84);
or(z124, t_1584, t_1585);
and(a125, f84, m122);
and(b125, m122, r74, n75, k74, h74);
not(t_1586, r120);
not(t_1587, w122);
or(c125, t_1586, t_1587);
and(d125, m122, r74, n75, k74);
and(e125, m122, r74, k74);
not(t_1588, s120);
not(t_1589, x122);
or(f125, t_1588, t_1589);
and(g125, m122, r74);
not(t_1590, k123);
not(t_1591, z112);
or(h125, t_1590, t_1591);
not(t_1592, d123);
not(t_1593, b113);
or(i125, t_1592, t_1593);
or(j125, a121, z122);
not(t_1594, e123);
not(t_1595, m113);
or(k125, t_1594, t_1595);
not(t_1596, b123);
not(t_1597, r113);
or(l125, t_1596, t_1597);
not(t_1598, c123);
not(t_1599, o108);
or(m125, t_1598, t_1599);
not(t_1600, g123);
not(t_1601, u113);
or(n125, t_1600, t_1601);
not(o125, m123);
not(t_1602, i121);
not(t_1603, n123);
or(p125, t_1602, t_1603);
not(t_1604, j121);
not(t_1605, o123);
or(q125, t_1604, t_1605);
not(t_1606, k121);
not(t_1607, p123);
or(r125, t_1606, t_1607);
not(t_1608, m121);
not(t_1609, q123);
or(s125, t_1608, t_1609);
not(t125, r123);
not(t_1610, v123);
not(t_1611, x101);
or(u125, t_1610, t_1611);
not(t_1612, w123);
not(t_1613, y101);
or(v125, t_1612, t_1613);
and(w125, n90, a124);
and(x125, a124, n79, k79, m79, h79);
and(y125, a124, n79, k79, m79);
not(t_1614, t121);
not(t_1615, x123);
or(z125, t_1614, t_1615);
not(t_1616, u121);
not(t_1617, y123);
or(a126, t_1616, t_1617);
and(b126, a124, n79, m79);
and(c126, a124, n79);
not(d126, z123);
buf(e126, a124);
not(t_1618, d124);
not(t_1619, v103);
or(f126, t_1618, t_1619);
not(t_1620, e124);
not(t_1621, w103);
or(g126, t_1620, t_1621);
not(t_1622, o125);
not(t_1623, n111);
or(h126, t_1622, t_1623);
not(t_1624, i122);
not(t_1625, i124);
or(i126, t_1624, t_1625);
not(j126, k124);
not(k126, l124);
not(t_1626, n122);
not(t_1627, m124);
or(l126, t_1626, t_1627);
not(t_1628, o122);
not(t_1629, n124);
or(m126, t_1628, t_1629);
or(n126, o124, d96);
not(t_1630, b106);
not(t_1631, r124);
or(o126, t_1630, t_1631);
not(t_1632, c106);
not(t_1633, t124);
or(p126, t_1632, t_1633);
or(q126, p124, q83, c83, p82, v37);
or(r126, q124, t83, e83, a38);
not(s126, r124);
or(t126, s124, s83, f38);
not(u126, t124);
or(v126, u124, k38);
not(t_1634, w96);
not(t_1635, r123);
or(w126, t_1634, t_1635);
not(t_1636, m49);
not(t_1637, x124);
or(x126, t_1636, t_1637);
not(t_1638, p49);
not(t_1639, w124);
or(y126, t_1638, t_1639);
not(z126, w124);
not(a127, x124);
and(b127, p106, z124);
or(c127, a125, a97);
and(d127, q106, y124);
not(t_1640, r106);
not(t_1641, c125);
or(e127, t_1640, t_1641);
not(t_1642, s106);
not(t_1643, f125);
or(f127, t_1642, t_1643);
or(g127, b125, j85, t84, q86, e39);
not(h127, c125);
or(i127, e125, l85, j39);
not(j127, f125);
or(k127, g125, o39);
not(t_1644, v97);
not(t_1645, l124);
or(l127, t_1644, t_1645);
not(t_1646, y122);
not(t_1647, h125);
or(m127, t_1646, t_1647);
not(t_1648, a123);
not(t_1649, i125);
or(n127, t_1648, t_1649);
not(t_1650, j125);
not(t_1651, p98);
or(o127, t_1650, t_1651);
or(p127, d125, m85, v84, d41);
not(t_1652, f123);
not(t_1653, k125);
or(q127, t_1652, t_1653);
not(t_1654, h123);
not(t_1655, l125);
or(r127, t_1654, t_1655);
not(t_1656, i123);
not(t_1657, m125);
or(s127, t_1656, t_1657);
not(t_1658, j123);
not(t_1659, n125);
or(t127, t_1658, t_1659);
not(t_1660, t123);
not(t_1661, u125);
or(u127, t_1660, t_1661);
not(t_1662, u123);
not(t_1663, v125);
or(v127, t_1662, t_1663);
or(w127, w125, o102);
or(x127, x125, q91, e91, v90, l46);
not(t_1664, c110);
not(t_1665, z125);
or(y127, t_1664, t_1665);
not(t_1666, d110);
not(t_1667, a126);
or(z127, t_1666, t_1667);
or(a128, y125, t91, g91, n46);
or(b128, b126, s91, p46);
not(c128, z125);
not(d128, a126);
or(e128, c126, r46);
not(t_1668, i103);
not(t_1669, e126);
or(f128, t_1668, t_1669);
not(g128, e126);
not(t_1670, b124);
not(t_1671, f126);
or(h128, t_1670, t_1671);
not(t_1672, c124);
not(t_1673, g126);
or(i128, t_1672, t_1673);
not(t_1674, h111);
not(t_1675, i126);
or(j128, t_1674, t_1675);
not(t_1676, h124);
not(t_1677, h126);
or(k128, t_1676, t_1677);
not(l128, i126);
and(m128, v124, j124, q127, t127);
and(n128, n126, o116);
and(o128, n126, r116);
not(p128, l126);
not(q128, m126);
and(r128, n126, t81);
and(s128, n126, t116);
not(t_1678, t95);
not(t_1679, l126);
or(t128, t_1678, t_1679);
not(t_1680, u95);
not(t_1681, m126);
or(u128, t_1680, t_1681);
not(v128, n126);
not(t_1682, e96);
not(t_1683, q126);
or(w128, t_1682, t_1683);
not(t_1684, s126);
not(t_1685, f96);
or(x128, t_1684, t_1685);
not(t_1686, u126);
not(t_1687, g96);
or(y128, t_1686, t_1687);
not(z128, q126);
not(t_1688, h96);
not(t_1689, r126);
or(a129, t_1688, t_1689);
not(b129, r126);
not(t_1690, p96);
not(t_1691, t126);
or(c129, t_1690, t_1691);
not(d129, t126);
not(t_1692, r96);
not(t_1693, v126);
or(e129, t_1692, t_1693);
not(f129, v126);
not(t_1694, t125);
not(t_1695, y83);
or(g129, t_1694, t_1695);
and(h129, b127, g49);
and(i129, c74, c127);
not(t_1696, a127);
not(t_1697, t38);
or(j129, t_1696, t_1697);
not(t_1698, z126);
not(t_1699, u38);
or(k129, t_1698, t_1699);
and(l129, c127, t49);
not(m129, b127);
not(n129, c127);
not(o129, d127);
not(t_1700, i97);
not(t_1701, g127);
or(p129, t_1700, t_1701);
not(t_1702, h127);
not(t_1703, j97);
or(q129, t_1702, t_1703);
not(t_1704, j127);
not(t_1705, k97);
or(r129, t_1704, t_1705);
not(s129, g127);
not(t_1706, l97);
not(t_1707, p127);
or(t129, t_1706, t_1707);
not(u129, i127);
not(t_1708, p97);
not(t_1709, k127);
or(v129, t_1708, t_1709);
not(w129, k127);
not(t_1710, k126);
not(t_1711, r85);
or(x129, t_1710, t_1711);
not(y129, p127);
not(t_1712, z98);
not(t_1713, i127);
or(z129, t_1712, t_1713);
and(a130, v113, o127);
and(b130, d127, s68);
and(c130, c127, b88);
and(d130, p125, q125, s127, m127);
and(e130, s125, r125, r127, n127);
and(f130, w78, o129);
and(g130, w127, q118);
not(h130, u127);
not(i130, v127);
and(j130, w127, u118);
not(t_1714, l102);
not(t_1715, u127);
or(k130, t_1714, t_1715);
not(t_1716, m102);
not(t_1717, v127);
or(l130, t_1716, t_1717);
and(m130, w127, j90);
and(n130, w127, x118);
not(o130, w127);
not(t_1718, t102);
not(t_1719, x127);
or(p130, t_1718, t_1719);
not(q130, x127);
not(t_1720, c128);
not(t_1721, u102);
or(r130, t_1720, t_1721);
not(t_1722, d128);
not(t_1723, v102);
or(s130, t_1722, t_1723);
not(t_1724, w102);
not(t_1725, a128);
or(t130, t_1724, t_1725);
not(u130, a128);
not(t_1726, d103);
not(t_1727, b128);
or(v130, t_1726, t_1727);
not(w130, b128);
not(t_1728, h103);
not(t_1729, e128);
or(x130, t_1728, t_1729);
not(y130, e128);
not(t_1730, g128);
not(t_1731, a92);
or(z130, t_1730, t_1731);
not(a131, h128);
not(b131, i128);
not(t_1732, j104);
not(t_1733, h128);
or(c131, t_1732, t_1733);
not(t_1734, k104);
not(t_1735, i128);
or(d131, t_1734, t_1735);
not(t_1736, l128);
not(t_1737, t104);
or(e131, t_1736, t_1737);
not(t_1738, f116);
not(t_1739, k128);
or(f131, t_1738, t_1739);
not(g131, k128);
and(h131, e130, m128, d130);
and(i131, y119, v128);
and(j131, d120, v128);
and(k131, a112, v128);
and(l131, c73, v128);
not(t_1740, p128);
not(t_1741, u81);
or(m131, t_1740, t_1741);
not(t_1742, q128);
not(t_1743, v81);
or(n131, t_1742, t_1743);
not(t_1744, z128);
not(t_1745, e82);
or(o131, t_1744, t_1745);
not(t_1746, o126);
not(t_1747, x128);
or(p131, t_1746, t_1747);
not(t_1748, p126);
not(t_1749, y128);
or(q131, t_1748, t_1749);
not(t_1750, b129);
not(t_1751, h82);
or(r131, t_1750, t_1751);
not(t_1752, d129);
not(t_1753, w82);
or(s131, t_1752, t_1753);
not(t_1754, f129);
not(t_1755, f83);
or(t131, t_1754, t_1755);
and(u131, a74, m129);
and(v131, h49, n129);
not(t_1756, x126);
not(t_1757, j129);
or(w131, t_1756, t_1757);
not(t_1758, y126);
not(t_1759, k129);
or(x131, t_1758, t_1759);
and(y131, x38, n129);
not(t_1760, s129);
not(t_1761, g84);
or(z131, t_1760, t_1761);
not(t_1762, e127);
not(t_1763, q129);
or(a132, t_1762, t_1763);
not(t_1764, f127);
not(t_1765, r129);
or(b132, t_1764, t_1765);
not(t_1766, y129);
not(t_1767, j84);
or(c132, t_1766, t_1767);
not(t_1768, w129);
not(t_1769, w84);
or(d132, t_1768, t_1769);
not(t_1770, u129);
not(t_1771, u86);
or(e132, t_1770, t_1771);
and(f132, a130, n108);
not(g132, a130);
and(h132, n77, n129);
and(i132, p121, o130);
and(j132, q121, o130);
and(k132, e115, o130);
not(t_1772, h130);
not(t_1773, h90);
or(l132, t_1772, t_1773);
not(t_1774, i130);
not(t_1775, i90);
or(m132, t_1774, t_1775);
and(n132, e79, o130);
not(t_1776, q130);
not(t_1777, o90);
or(o132, t_1776, t_1777);
not(t_1778, y127);
not(t_1779, r130);
or(p132, t_1778, t_1779);
not(t_1780, z127);
not(t_1781, s130);
or(q132, t_1780, t_1781);
not(t_1782, u130);
not(t_1783, r90);
or(r132, t_1782, t_1783);
not(t_1784, w130);
not(t_1785, d91);
or(s132, t_1784, t_1785);
not(t_1786, y130);
not(t_1787, p91);
or(t132, t_1786, t_1787);
not(t_1788, a131);
not(t_1789, m93);
or(u132, t_1788, t_1789);
not(t_1790, b131);
not(t_1791, n93);
or(v132, t_1790, t_1791);
not(t_1792, j128);
not(t_1793, e131);
or(w132, t_1792, t_1793);
not(t_1794, g131);
not(t_1795, i111);
or(x132, t_1794, t_1795);
not(t_1796, t128);
not(t_1797, m131);
or(y132, t_1796, t_1797);
not(t_1798, u128);
not(t_1799, n131);
or(z132, t_1798, t_1799);
not(a133, p131);
not(b133, q131);
not(t_1800, u96);
not(t_1801, p131);
or(c133, t_1800, t_1801);
not(t_1802, v96);
not(t_1803, q131);
or(d133, t_1802, t_1803);
or(e133, l129, y131);
and(f133, w131, z96, j126);
and(g133, x131, p106, j126);
and(h133, x131, p112, k124);
and(i133, w131, e117, k124);
not(j133, a132);
not(k133, b132);
not(t_1804, t97);
not(t_1805, a132);
or(l133, t_1804, t_1805);
not(t_1806, u97);
not(t_1807, b132);
or(m133, t_1806, t_1807);
and(n133, t18, s18, h131);
and(o133, u117, g132);
or(p133, c130, h132);
not(t_1808, k130);
not(t_1809, l132);
or(q133, t_1808, t_1809);
not(t_1810, l130);
not(t_1811, m132);
or(r133, t_1810, t_1811);
not(s133, p132);
not(t133, q132);
not(t_1812, j103);
not(t_1813, p132);
or(u133, t_1812, t_1813);
not(t_1814, k103);
not(t_1815, q132);
or(v133, t_1814, t_1815);
not(t_1816, c131);
not(t_1817, u132);
or(w133, t_1816, t_1817);
not(t_1818, d131);
not(t_1819, v132);
or(x133, t_1818, t_1819);
not(y133, w132);
not(t_1820, f131);
not(t_1821, x132);
or(z133, t_1820, t_1821);
not(t_1822, n95);
not(t_1823, z132);
or(a134, t_1822, t_1823);
not(t_1824, o95);
not(t_1825, y132);
or(b134, t_1824, t_1825);
not(c134, y132);
not(d134, z132);
not(t_1826, a133);
not(t_1827, u83);
or(e134, t_1826, t_1827);
not(t_1828, b133);
not(t_1829, v83);
or(f134, t_1828, t_1829);
or(g134, i133, h133, f133, g133);
not(t_1830, j133);
not(t_1831, n85);
or(h134, t_1830, t_1831);
not(t_1832, k133);
not(t_1833, o85);
or(i134, t_1832, t_1833);
not(t_1834, e114);
not(t_1835, w132);
or(j134, t_1834, t_1835);
not(t_1836, i102);
not(t_1837, r133);
or(k134, t_1836, t_1837);
not(t_1838, j102);
not(t_1839, q133);
or(l134, t_1838, t_1839);
not(m134, q133);
not(n134, r133);
not(t_1840, s133);
not(t_1841, b92);
or(o134, t_1840, t_1841);
not(t_1842, t133);
not(t_1843, c92);
or(p134, t_1842, t_1843);
not(t_1844, e104);
not(t_1845, x133);
or(q134, t_1844, t_1845);
not(t_1846, f104);
not(t_1847, w133);
or(r134, t_1846, t_1847);
not(s134, w133);
not(t134, x133);
not(u134, z133);
not(t_1848, d134);
not(t_1849, f81);
or(v134, t_1848, t_1849);
not(t_1850, c134);
not(t_1851, g81);
or(w134, t_1850, t_1851);
not(t_1852, c133);
not(t_1853, e134);
or(x134, t_1852, t_1853);
not(t_1854, d133);
not(t_1855, f134);
or(y134, t_1854, t_1855);
not(z134, g134);
not(t_1856, l133);
not(t_1857, h134);
or(a135, t_1856, t_1857);
not(t_1858, m133);
not(t_1859, i134);
or(b135, t_1858, t_1859);
not(t_1860, y133);
not(t_1861, a109);
or(c135, t_1860, t_1861);
not(t_1862, f114);
not(t_1863, z133);
or(d135, t_1862, t_1863);
not(t_1864, n134);
not(t_1865, w89);
or(e135, t_1864, t_1865);
not(t_1866, m134);
not(t_1867, x89);
or(f135, t_1866, t_1867);
not(t_1868, u133);
not(t_1869, o134);
or(g135, t_1868, t_1869);
not(t_1870, v133);
not(t_1871, p134);
or(h135, t_1870, t_1871);
not(t_1872, t134);
not(t_1873, y92);
or(i135, t_1872, t_1873);
not(t_1874, s134);
not(t_1875, z92);
or(j135, t_1874, t_1875);
not(t_1876, a134);
not(t_1877, v134);
or(k135, t_1876, t_1877);
not(t_1878, b134);
not(t_1879, w134);
or(l135, t_1878, t_1879);
not(t_1880, s96);
not(t_1881, y134);
or(m135, t_1880, t_1881);
not(t_1882, t96);
not(t_1883, x134);
or(n135, t_1882, t_1883);
not(o135, x134);
not(p135, y134);
not(t_1884, r97);
not(t_1885, b135);
or(q135, t_1884, t_1885);
not(t_1886, s97);
not(t_1887, a135);
or(r135, t_1886, t_1887);
not(s135, a135);
not(t135, b135);
not(t_1888, j134);
not(t_1889, c135);
or(u135, t_1888, t_1889);
not(t_1890, u134);
not(t_1891, b109);
or(v135, t_1890, t_1891);
not(t_1892, k134);
not(t_1893, e135);
or(w135, t_1892, t_1893);
not(t_1894, l134);
not(t_1895, f135);
or(x135, t_1894, t_1895);
not(t_1896, f103);
not(t_1897, h135);
or(y135, t_1896, t_1897);
not(t_1898, g103);
not(t_1899, g135);
or(z135, t_1898, t_1899);
not(a136, g135);
not(b136, h135);
not(t_1900, q134);
not(t_1901, i135);
or(c136, t_1900, t_1901);
not(t_1902, r134);
not(t_1903, j135);
or(d136, t_1902, t_1903);
not(t_1904, f105);
not(t_1905, u135);
or(e136, t_1904, t_1905);
not(t_1906, u94);
not(t_1907, l135);
or(f136, t_1906, t_1907);
not(t_1908, v94);
not(t_1909, k135);
or(g136, t_1908, t_1909);
not(h136, k135);
not(i136, l135);
not(t_1910, p135);
not(t_1911, g83);
or(j136, t_1910, t_1911);
not(t_1912, o135);
not(t_1913, h83);
or(k136, t_1912, t_1913);
not(t_1914, t135);
not(t_1915, z84);
or(l136, t_1914, t_1915);
not(t_1916, s135);
not(t_1917, b85);
or(m136, t_1916, t_1917);
not(n136, u135);
not(t_1918, d135);
not(t_1919, v135);
or(o136, t_1918, t_1919);
not(t_1920, q101);
not(t_1921, x135);
or(p136, t_1920, t_1921);
not(t_1922, r101);
not(t_1923, w135);
or(q136, t_1922, t_1923);
not(r136, w135);
not(s136, x135);
not(t_1924, b136);
not(t_1925, m91);
or(t136, t_1924, t_1925);
not(t_1926, a136);
not(t_1927, n91);
or(u136, t_1926, t_1927);
not(t_1928, o103);
not(t_1929, d136);
or(v136, t_1928, t_1929);
not(t_1930, p103);
not(t_1931, c136);
or(w136, t_1930, t_1931);
not(x136, c136);
not(y136, d136);
not(t_1932, e105);
not(t_1933, o136);
or(z136, t_1932, t_1933);
not(t_1934, n136);
not(t_1935, o94);
or(a137, t_1934, t_1935);
not(t_1936, i136);
not(t_1937, i80);
or(b137, t_1936, t_1937);
not(t_1938, h136);
not(t_1939, j80);
or(c137, t_1938, t_1939);
not(t_1940, m135);
not(t_1941, j136);
or(d137, t_1940, t_1941);
not(t_1942, n135);
not(t_1943, k136);
or(e137, t_1942, t_1943);
not(t_1944, q135);
not(t_1945, l136);
or(f137, t_1944, t_1945);
not(t_1946, r135);
not(t_1947, m136);
or(g137, t_1946, t_1947);
not(h137, o136);
not(t_1948, s136);
not(t_1949, z88);
or(i137, t_1948, t_1949);
not(t_1950, r136);
not(t_1951, a89);
or(j137, t_1950, t_1951);
not(t_1952, y135);
not(t_1953, t136);
or(k137, t_1952, t_1953);
not(t_1954, z135);
not(t_1955, u136);
or(l137, t_1954, t_1955);
not(t_1956, y136);
not(t_1957, e92);
or(m137, t_1956, t_1957);
not(t_1958, x136);
not(t_1959, f92);
or(n137, t_1958, t_1959);
not(t_1960, h137);
not(t_1961, n94);
or(o137, t_1960, t_1961);
not(t_1962, e136);
not(t_1963, a137);
or(p137, t_1962, t_1963);
not(t_1964, f136);
not(t_1965, b137);
or(q137, t_1964, t_1965);
not(t_1966, g136);
not(t_1967, c137);
or(r137, t_1966, t_1967);
not(t_1968, a96);
not(t_1969, e137);
or(s137, t_1968, t_1969);
not(t_1970, b96);
not(t_1971, d137);
or(t137, t_1970, t_1971);
not(u137, d137);
not(v137, e137);
not(t_1972, f97);
not(t_1973, g137);
or(w137, t_1972, t_1973);
not(t_1974, g97);
not(t_1975, f137);
or(x137, t_1974, t_1975);
not(y137, f137);
not(z137, g137);
not(t_1976, p136);
not(t_1977, i137);
or(a138, t_1976, t_1977);
not(t_1978, q136);
not(t_1979, j137);
or(b138, t_1978, t_1979);
not(t_1980, q102);
not(t_1981, l137);
or(c138, t_1980, t_1981);
not(t_1982, r102);
not(t_1983, k137);
or(d138, t_1982, t_1983);
not(e138, k137);
not(f138, l137);
not(t_1984, v136);
not(t_1985, m137);
or(g138, t_1984, t_1985);
not(t_1986, w136);
not(t_1987, n137);
or(h138, t_1986, t_1987);
not(t_1988, q104);
not(t_1989, p137);
or(i138, t_1988, t_1989);
not(t_1990, z136);
not(t_1991, o137);
or(j138, t_1990, t_1991);
not(k138, p137);
not(l138, q137);
not(m138, r137);
not(t_1992, h95);
not(t_1993, r137);
or(n138, t_1992, t_1993);
not(t_1994, i95);
not(t_1995, q137);
or(o138, t_1994, t_1995);
not(t_1996, v137);
not(t_1997, a82);
or(p138, t_1996, t_1997);
not(t_1998, u137);
not(t_1999, b82);
or(q138, t_1998, t_1999);
not(t_2000, z137);
not(t_2001, c84);
or(r138, t_2000, t_2001);
not(t_2002, y137);
not(t_2003, d84);
or(s138, t_2002, t_2003);
not(t138, a138);
not(u138, b138);
not(t_2004, b102);
not(t_2005, b138);
or(v138, t_2004, t_2005);
not(t_2006, c102);
not(t_2007, a138);
or(w138, t_2006, t_2007);
not(t_2008, f138);
not(t_2009, k90);
or(x138, t_2008, t_2009);
not(t_2010, e138);
not(t_2011, l90);
or(y138, t_2010, t_2011);
not(z138, g138);
not(a139, h138);
not(t_2012, z103);
not(t_2013, h138);
or(b139, t_2012, t_2013);
not(t_2014, a104);
not(t_2015, g138);
or(c139, t_2014, t_2015);
not(t_2016, k138);
not(t_2017, q93);
or(d139, t_2016, t_2017);
not(t_2018, r104);
not(t_2019, j138);
or(e139, t_2018, t_2019);
not(f139, j138);
not(t_2020, m138);
not(t_2021, t80);
or(g139, t_2020, t_2021);
not(t_2022, l138);
not(t_2023, v80);
or(h139, t_2022, t_2023);
not(t_2024, s137);
not(t_2025, p138);
or(i139, t_2024, t_2025);
not(t_2026, t137);
not(t_2027, q138);
or(j139, t_2026, t_2027);
not(t_2028, w137);
not(t_2029, r138);
or(k139, t_2028, t_2029);
not(t_2030, x137);
not(t_2031, s138);
or(l139, t_2030, t_2031);
not(t_2032, u138);
not(t_2033, j89);
or(m139, t_2032, t_2033);
not(t_2034, t138);
not(t_2035, l89);
or(n139, t_2034, t_2035);
not(t_2036, c138);
not(t_2037, x138);
or(o139, t_2036, t_2037);
not(t_2038, d138);
not(t_2039, y138);
or(p139, t_2038, t_2039);
not(t_2040, a139);
not(t_2041, o92);
or(q139, t_2040, t_2041);
not(t_2042, z138);
not(t_2043, q92);
or(r139, t_2042, t_2043);
not(t_2044, i138);
not(t_2045, d139);
or(s139, t_2044, t_2045);
not(t_2046, f139);
not(t_2047, r93);
or(t139, t_2046, t_2047);
not(t_2048, n138);
not(t_2049, g139);
or(u139, t_2048, t_2049);
not(t_2050, o138);
not(t_2051, h139);
or(v139, t_2050, t_2051);
not(w139, i139);
not(x139, j139);
not(t_2052, n96);
not(t_2053, i139);
or(y139, t_2052, t_2053);
not(t_2054, o96);
not(t_2055, j139);
or(z139, t_2054, t_2055);
not(a140, k139);
not(b140, l139);
not(t_2056, x98);
not(t_2057, k139);
or(c140, t_2056, t_2057);
not(t_2058, y98);
not(t_2059, l139);
or(d140, t_2058, t_2059);
not(t_2060, v138);
not(t_2061, m139);
or(e140, t_2060, t_2061);
not(t_2062, w138);
not(t_2063, n139);
or(f140, t_2062, t_2063);
not(g140, o139);
not(h140, p139);
not(t_2064, b103);
not(t_2065, o139);
or(i140, t_2064, t_2065);
not(t_2066, c103);
not(t_2067, p139);
or(j140, t_2066, t_2067);
not(t_2068, b139);
not(t_2069, q139);
or(k140, t_2068, t_2069);
not(t_2070, c139);
not(t_2071, r139);
or(l140, t_2070, t_2071);
not(m140, s139);
not(t_2072, e139);
not(t_2073, t139);
or(n140, t_2072, t_2073);
not(t_2074, a105);
not(t_2075, s139);
or(o140, t_2074, t_2075);
and(p140, u139, z95, s123);
and(q140, v139, a106, s123);
and(r140, v139, e112, o121);
and(s140, u139, w116, o121);
not(t_2076, w139);
not(t_2077, t82);
or(t140, t_2076, t_2077);
not(t_2078, x139);
not(t_2079, u82);
or(u140, t_2078, t_2079);
not(t_2080, a140);
not(t_2081, s86);
or(v140, t_2080, t_2081);
not(t_2082, b140);
not(t_2083, t86);
or(w140, t_2082, t_2083);
and(x140, l140, c116, n13);
and(y140, k140, m119, n13);
and(z140, l140, e111, e16);
and(a141, k140, n104, e16);
and(b141, e140, p102, d126);
and(c141, f140, b110, d126);
and(d141, f140, i115, z123);
and(e141, e140, y118, z123);
not(t_2084, g140);
not(t_2085, a91);
or(f141, t_2084, t_2085);
not(t_2086, h140);
not(t_2087, b91);
or(g141, t_2086, t_2087);
not(h141, n140);
not(t_2088, m140);
not(t_2089, d94);
or(i141, t_2088, t_2089);
not(t_2090, b105);
not(t_2091, n140);
or(j141, t_2090, t_2091);
or(k141, s140, r140, p140, q140);
not(t_2092, y139);
not(t_2093, t140);
or(l141, t_2092, t_2093);
not(t_2094, z139);
not(t_2095, u140);
or(m141, t_2094, t_2095);
not(t_2096, c140);
not(t_2097, v140);
or(n141, t_2096, t_2097);
not(t_2098, d140);
not(t_2099, w140);
or(o141, t_2098, t_2099);
or(p141, y140, x140, a141, z140);
or(q141, e141, d141, b141, c141);
not(t_2100, i140);
not(t_2101, f141);
or(r141, t_2100, t_2101);
not(t_2102, j140);
not(t_2103, g141);
or(s141, t_2102, t_2103);
not(t_2104, o140);
not(t_2105, i141);
or(t141, t_2104, t_2105);
not(t_2106, h141);
not(t_2107, e94);
or(u141, t_2106, t_2107);
not(v141, k141);
not(t_2108, i96);
not(t_2109, l141);
or(w141, t_2108, t_2109);
not(t_2110, j96);
not(t_2111, m141);
or(x141, t_2110, t_2111);
not(y141, l141);
not(z141, m141);
not(t_2112, m97);
not(t_2113, n141);
or(a142, t_2112, t_2113);
not(t_2114, n97);
not(t_2115, o141);
or(b142, t_2114, t_2115);
not(c142, n141);
not(d142, o141);
not(e142, p141);
not(f142, q141);
not(t_2116, x102);
not(t_2117, r141);
or(g142, t_2116, t_2117);
not(t_2118, y102);
not(t_2119, s141);
or(h142, t_2118, t_2119);
not(i142, r141);
not(j142, s141);
not(t_2120, u104);
not(t_2121, t141);
or(k142, t_2120, t_2121);
not(l142, t141);
not(t_2122, j141);
not(t_2123, u141);
or(m142, t_2122, t_2123);
not(t_2124, y141);
not(t_2125, i82);
or(n142, t_2124, t_2125);
not(t_2126, z141);
not(t_2127, k82);
or(o142, t_2126, t_2127);
not(t_2128, c142);
not(t_2129, k84);
or(p142, t_2128, t_2129);
not(t_2130, d142);
not(t_2131, m84);
or(q142, t_2130, t_2131);
not(t_2132, i142);
not(t_2133, s90);
or(r142, t_2132, t_2133);
not(t_2134, j142);
not(t_2135, u90);
or(s142, t_2134, t_2135);
not(t_2136, l142);
not(t_2137, u93);
or(t142, t_2136, t_2137);
not(t_2138, w104);
not(t_2139, m142);
or(u142, t_2138, t_2139);
not(v142, m142);
not(t_2140, w141);
not(t_2141, n142);
or(w142, t_2140, t_2141);
not(t_2142, x141);
not(t_2143, o142);
or(x142, t_2142, t_2143);
not(t_2144, a142);
not(t_2145, p142);
or(y142, t_2144, t_2145);
not(t_2146, b142);
not(t_2147, q142);
or(z142, t_2146, t_2147);
and(a143, o121, x142);
not(t_2148, g142);
not(t_2149, r142);
or(b143, t_2148, t_2149);
not(t_2150, h142);
not(t_2151, s142);
or(c143, t_2150, t_2151);
not(t_2152, k142);
not(t_2153, t142);
or(d143, t_2152, t_2153);
not(t_2154, v142);
not(t_2155, v93);
or(e143, t_2154, t_2155);
and(f143, k124, z142);
not(g143, w142);
not(h143, y142);
and(i143, g143, s123);
not(j143, b143);
and(k143, z123, c143);
not(l143, d143);
not(t_2156, u142);
not(t_2157, e143);
or(m143, t_2156, t_2157);
and(n143, h143, j126);
and(o143, n13, m143);
and(p143, l143, e16);
or(q143, a143, i143);
and(r143, j143, d126);
or(s143, f143, n143);
or(t143, o143, p143);
not(u143, q143);
or(v143, k143, r143);
not(w143, s143);
not(t_2158, v141);
not(t_2159, q143);
or(x143, t_2158, t_2159);
not(t_2160, z134);
not(t_2161, s143);
or(y143, t_2160, t_2161);
not(t_2162, e142);
not(t_2163, t143);
or(z143, t_2162, t_2163);
not(a144, t143);
not(t_2164, f142);
not(t_2165, v143);
or(b144, t_2164, t_2165);
not(c144, v143);
not(t_2166, u143);
not(t_2167, k141);
or(d144, t_2166, t_2167);
not(t_2168, w143);
not(t_2169, g134);
or(e144, t_2168, t_2169);
not(t_2170, a144);
not(t_2171, p141);
or(f144, t_2170, t_2171);
not(t_2172, c144);
not(t_2173, q141);
or(g144, t_2172, t_2173);
not(t_2174, d144);
not(t_2175, x143);
or(h144, t_2174, t_2175);
not(t_2176, e144);
not(t_2177, y143);
or(i144, t_2176, t_2177);
not(t_2178, f144);
not(t_2179, z143);
or(j144, t_2178, t_2179);
not(t_2180, g144);
not(t_2181, b144);
or(k144, t_2180, t_2181);
buf(z6, i5);
buf(a7, a);
buf(b7, a);
buf(c7, l5);
buf(d7, n5);
buf(e7, o5);
buf(f7, p5);
buf(g7, q5);
buf(h7, r5);
buf(i7, t5);
buf(j7, v5);
buf(k7, w5);
buf(l7, x5);
buf(m7, y5);
buf(n7, z5);
buf(o7, a6);
buf(p7, b6);
buf(q7, c6);
buf(r7, d6);
buf(s7, e6);
buf(t7, f6);
buf(u7, g6);
buf(v7, h6);
buf(w7, i6);
buf(x7, j6);
buf(y7, k6);
buf(z7, l6);
buf(a8, m6);
buf(b8, n6);
buf(c8, p6);
buf(d8, q6);
buf(e8, r6);
buf(f8, s6);
buf(g8, t6);
buf(h8, u6);
buf(i8, v6);
buf(j8, w6);
buf(l8, m5);
buf(m8, u5);
buf(n8, o6);
buf(n10, p133);
buf(o10, p133);
buf(p10, e133);
buf(q10, e133);
endmodule
module top;
	parameter in_width = 207,
		patterns = 5000,
		step = 1;
	reg [1:in_width] in_mem[1:patterns];
	integer index;

	wire i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,
		i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,
		i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,
		i30,i31,i32,i33,i34,i35,i36,i37,i38,i39,
		i40,i41,i42,i43,i44,i45,i46,i47,i48,i49,
		i50,i51,i52,i53,i54,i55,i56,i57,i58,i59,
		i60,i61,i62,i63,i64,i65,i66,i67,i68,i69,
		i70,i71,i72,i73,i74,i75,i76,i77,i78,i79,
		i80,i81,i82,i83,i84,i85,i86,i87,i88,i89,
		i90,i91,i92,i93,i94,i95,i96,i97,i98,i99,
		i100,i101,i102,i103,i104,i105,i106,i107,i108,i109,
		i110,i111,i112,i113,i114,i115,i116,i117,i118,i119,
		i120,i121,i122,i123,i124,i125,i126,i127,i128,i129,
		i130,i131,i132,i133,i134,i135,i136,i137,i138,i139,
		i140,i141,i142,i143,i144,i145,i146,i147,i148,i149,
		i150,i151,i152,i153,i154,i155,i156,i157,i158,i159,
		i160,i161,i162,i163,i164,i165,i166,i167,i168,i169,
		i170,i171,i172,i173,i174,i175,i176,i177,i178,i179,
		i180,i181,i182,i183,i184,i185,i186,i187,i188,i189,
		i190,i191,i192,i193,i194,i195,i196,i197,i198,i199,
		i200,i201,i202,i203,i204,i205,i206;

	assign {i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,
		i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,
		i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,
		i30,i31,i32,i33,i34,i35,i36,i37,i38,i39,
		i40,i41,i42,i43,i44,i45,i46,i47,i48,i49,
		i50,i51,i52,i53,i54,i55,i56,i57,i58,i59,
		i60,i61,i62,i63,i64,i65,i66,i67,i68,i69,
		i70,i71,i72,i73,i74,i75,i76,i77,i78,i79,
		i80,i81,i82,i83,i84,i85,i86,i87,i88,i89,
		i90,i91,i92,i93,i94,i95,i96,i97,i98,i99,
		i100,i101,i102,i103,i104,i105,i106,i107,i108,i109,
		i110,i111,i112,i113,i114,i115,i116,i117,i118,i119,
		i120,i121,i122,i123,i124,i125,i126,i127,i128,i129,
		i130,i131,i132,i133,i134,i135,i136,i137,i138,i139,
		i140,i141,i142,i143,i144,i145,i146,i147,i148,i149,
		i150,i151,i152,i153,i154,i155,i156,i157,i158,i159,
		i160,i161,i162,i163,i164,i165,i166,i167,i168,i169,
		i170,i171,i172,i173,i174,i175,i176,i177,i178,i179,
		i180,i181,i182,i183,i184,i185,i186,i187,i188,i189,
		i190,i191,i192,i193,i194,i195,i196,i197,i198,i199,
		i200,i201,i202,i203,i204,i205,i206} = 
		$getpattern(in_mem[index]);

	initial $monitor($time,,o0,o1,o2,o3,o4,o5,o6,o7,o8,o9,
		o10,o11,o12,o13,o14,o15,o16,o17,o18,o19,
		o20,o21,o22,o23,o24,o25,o26,o27,o28,o29,
		o30,o31,o32,o33,o34,o35,o36,o37,o38,o39,
		o40,o41,o42,o43,o44,o45,o46,o47,o48,o49,
		o50,o51,o52,o53,o54,o55,o56,o57,o58,o59,
		o60,o61,o62,o63,o64,o65,o66,o67,o68,o69,
		o70,o71,o72,o73,o74,o75,o76,o77,o78,o79,
		o80,o81,o82,o83,o84,o85,o86,o87,o88,o89,
		o90,o91,o92,o93,o94,o95,o96,o97,o98,o99,
		o100,o101,o102,o103,o104,o105,o106,o107);
	initial
		begin
			$readmemb("patt.mem", in_mem);
			for(index = 1; index <= patterns; index = index + 1)
				#step;
		end

	foobar cct(o0,o1,o2,o3,o4,o5,o6,o7,o8,o9,
		o10,o11,o12,o13,o14,o15,o16,o17,o18,o19,
		o20,o21,o22,o23,o24,o25,o26,o27,o28,o29,
		o30,o31,o32,o33,o34,o35,o36,o37,o38,o39,
		o40,o41,o42,o43,o44,o45,o46,o47,o48,o49,
		o50,o51,o52,o53,o54,o55,o56,o57,o58,o59,
		o60,o61,o62,o63,o64,o65,o66,o67,o68,o69,
		o70,o71,o72,o73,o74,o75,o76,o77,o78,o79,
		o80,o81,o82,o83,o84,o85,o86,o87,o88,o89,
		o90,o91,o92,o93,o94,o95,o96,o97,o98,o99,
		o100,o101,o102,o103,o104,o105,o106,o107,i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,
		i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,
		i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,
		i30,i31,i32,i33,i34,i35,i36,i37,i38,i39,
		i40,i41,i42,i43,i44,i45,i46,i47,i48,i49,
		i50,i51,i52,i53,i54,i55,i56,i57,i58,i59,
		i60,i61,i62,i63,i64,i65,i66,i67,i68,i69,
		i70,i71,i72,i73,i74,i75,i76,i77,i78,i79,
		i80,i81,i82,i83,i84,i85,i86,i87,i88,i89,
		i90,i91,i92,i93,i94,i95,i96,i97,i98,i99,
		i100,i101,i102,i103,i104,i105,i106,i107,i108,i109,
		i110,i111,i112,i113,i114,i115,i116,i117,i118,i119,
		i120,i121,i122,i123,i124,i125,i126,i127,i128,i129,
		i130,i131,i132,i133,i134,i135,i136,i137,i138,i139,
		i140,i141,i142,i143,i144,i145,i146,i147,i148,i149,
		i150,i151,i152,i153,i154,i155,i156,i157,i158,i159,
		i160,i161,i162,i163,i164,i165,i166,i167,i168,i169,
		i170,i171,i172,i173,i174,i175,i176,i177,i178,i179,
		i180,i181,i182,i183,i184,i185,i186,i187,i188,i189,
		i190,i191,i192,i193,i194,i195,i196,i197,i198,i199,
		i200,i201,i202,i203,i204,i205,i206);
endmodule
