// IWLS benchmark module "apex6" printed on Wed May 29 16:03:29 2002
module apex6(PSRW, VFIN, PFIN, INFIN, VYBB0, VYBB1, VZZZE, PYBB0, PYBB1, PYBB2, PYBB3, PYBB4, PYBB5, PYBB6, PYBB7, PYBB8, PZZZE, INYBB0, INYBB1, INYBB2, INYBB3, INYBB4, INYBB5, INYBB6, INYBB7, INYBB8, INZZZE, MMERR, ESRSUM, CBT0, CBT1, CBT2, SLAD0, SLAD1, SLAD2, SLAD3, PSYNC, RPTEN, ICLR, STW_N, P1ZZZ0, P1ZZZ1, P1ZZZ2, P1ZZZ3, P1ZZZ4, P1ZZZ5, P1ZZZ6, P1ZZZ7, P2ZZZ0, P2ZZZ1, P2ZZZ2, P2ZZZ3, P2ZZZ4, P2ZZZ5, P2ZZZ6, P2ZZZ7, I1ZZZ0, I1ZZZ1, I1ZZZ2, I1ZZZ3, I1ZZZ4, I1ZZZ5, I1ZZZ6, I1ZZZ7, I2ZZZ0, I2ZZZ1, I2ZZZ2, I2ZZZ3, I2ZZZ4, I2ZZZ5, I2ZZZ6, I2ZZZ7, TXMESS_N, RYZ, COMPPAR, RPTWIN, XZFR0, XZFR1, XZFS, RXZ0, RXZ1, OFS2, OFS1, A, B, C, QPR0, QPR1, QPR2, QPR3, QPR4, AXZ0, AXZ1, V1ZZZ0, V1ZZZ1, V1ZZZ2, V1ZZZ3, V1ZZZ4, V1ZZZ5, V1ZZZ6, V1ZZZ7, V2ZZZ0, V2ZZZ1, V2ZZZ2, V2ZZZ3, V2ZZZ4, V2ZZZ5, V2ZZZ6, V2ZZZ7, TXWRD0, TXWRD1, TXWRD2, TXWRD3, TXWRD4, TXWRD5, TXWRD6, TXWRD7, TXWRD8, TXWRD9, TXWRD10, TXWRD11, TXWRD12, TXWRD13, TXWRD14, TXWRD15, XZ320, XZ321, XZ322, XZ323, XZ324, XZ160_N, XZ161, XZ162, XZ163, ENWIN, SBUFF, STW_F, TD_P, FSESR_P, P1ZZZ0_P, P1ZZZ1_P, P1ZZZ2_P, P1ZZZ3_P, P1ZZZ4_P, P1ZZZ5_P, P1ZZZ6_P, P1ZZZ7_P, P2ZZZ0_P, P2ZZZ1_P, P2ZZZ2_P, P2ZZZ3_P, P2ZZZ4_P, P2ZZZ5_P, P2ZZZ6_P, P2ZZZ7_P, I1ZZZ0_P, I1ZZZ1_P, I1ZZZ2_P, I1ZZZ3_P, I1ZZZ4_P, I1ZZZ5_P, I1ZZZ6_P, I1ZZZ7_P, I2ZZZ0_P, I2ZZZ1_P, I2ZZZ2_P, I2ZZZ3_P, I2ZZZ4_P, I2ZZZ5_P, I2ZZZ6_P, I2ZZZ7_P, TXMESS_F, RYZ_P, COMPPAR_P, RPTWIN_P, XZFR0_P, XZFR1_P, XZFS_P, RXZ0_P, RXZ1_P, OFS2_P, OFS1_P, A_P, B_P, C_P, QPR0_P, QPR1_P, QPR2_P, QPR3_P, QPR4_P, AXZ0_P, AXZ1_P, V1ZZZ0_P, V1ZZZ1_P, V1ZZZ2_P, V1ZZZ3_P, V1ZZZ4_P, V1ZZZ5_P, V1ZZZ6_P, V1ZZZ7_P, V2ZZZ0_P, V2ZZZ1_P, V2ZZZ2_P, V2ZZZ3_P, V2ZZZ4_P, V2ZZZ5_P, V2ZZZ6_P, V2ZZZ7_P, TXWRD0_P, TXWRD1_P, TXWRD2_P, TXWRD3_P, TXWRD4_P, TXWRD5_P, TXWRD6_P, TXWRD7_P, TXWRD8_P, TXWRD9_P, TXWRD10_P, TXWRD11_P, TXWRD12_P, TXWRD13_P, TXWRD14_P, TXWRD15_P, XZ320_P, XZ321_P, XZ322_P, XZ323_P, XZ324_P, XZ160_F, XZ161_P, XZ162_P, XZ163_P, ENWIN_P);
input
  A,
  B,
  C,
  STW_N,
  QPR0,
  QPR1,
  QPR2,
  QPR3,
  QPR4,
  ENWIN,
  INZZZE,
  XZFR0,
  XZFR1,
  VZZZE,
  RXZ0,
  RXZ1,
  INFIN,
  V2ZZZ0,
  V2ZZZ1,
  V2ZZZ2,
  V2ZZZ3,
  V2ZZZ4,
  V2ZZZ5,
  V2ZZZ6,
  V2ZZZ7,
  XZ161,
  XZ162,
  XZ163,
  I2ZZZ0,
  I2ZZZ1,
  I2ZZZ2,
  I2ZZZ3,
  I2ZZZ4,
  I2ZZZ5,
  I2ZZZ6,
  XZ160_N,
  I2ZZZ7,
  TXMESS_N,
  PZZZE,
  RYZ,
  AXZ0,
  AXZ1,
  COMPPAR,
  MMERR,
  V1ZZZ0,
  PSRW,
  V1ZZZ1,
  V1ZZZ2,
  V1ZZZ3,
  V1ZZZ4,
  V1ZZZ5,
  V1ZZZ6,
  V1ZZZ7,
  I1ZZZ0,
  I1ZZZ1,
  I1ZZZ2,
  I1ZZZ3,
  I1ZZZ4,
  I1ZZZ5,
  I1ZZZ6,
  I1ZZZ7,
  RPTEN,
  XZ320,
  XZ321,
  XZ322,
  XZ323,
  XZ324,
  CBT0,
  CBT1,
  CBT2,
  ESRSUM,
  SLAD0,
  SLAD1,
  SLAD2,
  SLAD3,
  XZFS,
  RPTWIN,
  PFIN,
  PSYNC,
  OFS1,
  OFS2,
  P2ZZZ0,
  P2ZZZ1,
  P2ZZZ2,
  P2ZZZ3,
  P2ZZZ4,
  TXWRD0,
  P2ZZZ5,
  TXWRD1,
  P2ZZZ6,
  TXWRD2,
  P2ZZZ7,
  TXWRD3,
  TXWRD4,
  TXWRD5,
  TXWRD6,
  TXWRD7,
  TXWRD8,
  TXWRD9,
  INYBB0,
  INYBB1,
  INYBB2,
  INYBB3,
  INYBB4,
  INYBB5,
  INYBB6,
  INYBB7,
  INYBB8,
  VYBB0,
  VYBB1,
  TXWRD10,
  TXWRD11,
  TXWRD12,
  TXWRD13,
  TXWRD14,
  TXWRD15,
  PYBB0,
  PYBB1,
  PYBB2,
  PYBB3,
  PYBB4,
  PYBB5,
  PYBB6,
  PYBB7,
  PYBB8,
  ICLR,
  P1ZZZ0,
  P1ZZZ1,
  P1ZZZ2,
  P1ZZZ3,
  P1ZZZ4,
  P1ZZZ5,
  P1ZZZ6,
  P1ZZZ7,
  VFIN;
output
  V2ZZZ2_P,
  QPR3_P,
  XZ323_P,
  P1ZZZ4_P,
  I1ZZZ3_P,
  TXWRD5_P,
  STW_F,
  TXWRD13_P,
  V1ZZZ4_P,
  P2ZZZ1_P,
  I2ZZZ2_P,
  TXWRD0_P,
  A_P,
  V2ZZZ1_P,
  TXWRD8_P,
  QPR4_P,
  XZ324_P,
  P1ZZZ3_P,
  I1ZZZ4_P,
  V1ZZZ3_P,
  COMPPAR_P,
  XZFS_P,
  P2ZZZ4_P,
  I2ZZZ3_P,
  XZ160_F,
  B_P,
  TXMESS_F,
  TXWRD7_P,
  P1ZZZ6_P,
  V2ZZZ4_P,
  I1ZZZ5_P,
  TXWRD15_P,
  V1ZZZ6_P,
  XZ161_P,
  RPTWIN_P,
  P2ZZZ3_P,
  AXZ0_P,
  I2ZZZ4_P,
  TXWRD2_P,
  C_P,
  P1ZZZ5_P,
  V2ZZZ3_P,
  I1ZZZ6_P,
  FSESR_P,
  V1ZZZ5_P,
  XZ162_P,
  TXWRD10_P,
  P1ZZZ0_P,
  OFS1_P,
  P2ZZZ6_P,
  AXZ1_P,
  I2ZZZ5_P,
  TXWRD1_P,
  I1ZZZ7_P,
  TXWRD9_P,
  ENWIN_P,
  V1ZZZ0_P,
  V2ZZZ6_P,
  XZ163_P,
  OFS2_P,
  P2ZZZ5_P,
  I1ZZZ0_P,
  I2ZZZ6_P,
  QPR0_P,
  XZ320_P,
  P1ZZZ7_P,
  TXWRD4_P,
  RXZ0_P,
  V2ZZZ5_P,
  SBUFF,
  V1ZZZ7_P,
  P2ZZZ0_P,
  TXWRD12_P,
  I2ZZZ7_P,
  P1ZZZ2_P,
  V2ZZZ0_P,
  I1ZZZ1_P,
  QPR1_P,
  XZ321_P,
  TXWRD3_P,
  RXZ1_P,
  V1ZZZ2_P,
  XZFR0_P,
  TD_P,
  I2ZZZ0_P,
  P2ZZZ7_P,
  TXWRD11_P,
  P1ZZZ1_P,
  I1ZZZ2_P,
  RYZ_P,
  QPR2_P,
  XZ322_P,
  V2ZZZ7_P,
  TXWRD6_P,
  V1ZZZ1_P,
  XZFR1_P,
  TXWRD14_P,
  P2ZZZ2_P,
  I2ZZZ1_P;
wire
  \[60] ,
  MIS16871,
  MIS16873,
  MIS16879,
  \[61] ,
  \[62] ,
  MIS16891,
  MIS16893,
  MIS16895,
  \[63] ,
  \[64] ,
  \[65] ,
  \[66] ,
  \[67] ,
  MIS16701,
  MIS16706,
  \[68] ,
  MIS11154,
  \[69] ,
  MIS16722,
  MIS16724,
  MIS16726,
  MIS16728,
  MIS16710,
  MIS16712,
  MIS16716,
  MIS16719,
  MIS16740,
  MIS16742,
  MIS16746,
  MIS16748,
  \[0] ,
  MIS16730,
  MIS16732,
  MIS16734,
  MIS16736,
  \[1] ,
  MIS16760,
  MIS16762,
  MIS16765,
  MIS16767,
  \[2] ,
  MIS16750,
  MIS8768,
  MIS16752,
  MIS16754,
  MIS16758,
  \[3] ,
  MIS8027,
  MIS16780,
  MIS16786,
  MIS16788,
  \[4] ,
  \[70] ,
  MIS16778,
  \[5] ,
  \[71] ,
  \[6] ,
  \[72] ,
  MIS16790,
  MIS16792,
  \[7] ,
  \[73] ,
  \[8] ,
  \[74] ,
  \[9] ,
  \[75] ,
  \[76] ,
  \[77] ,
  \[78] ,
  \[79] ,
  MIS12425,
  \[80] ,
  \[81] ,
  MIS9061,
  \[82] ,
  \[83] ,
  MIS15964,
  \[84] ,
  MIS9071,
  \[85] ,
  \[86] ,
  \[87] ,
  \[88] ,
  \[89] ,
  \[10] ,
  \[11] ,
  \[12] ,
  \[13] ,
  \[90] ,
  \[14] ,
  \[91] ,
  \[15] ,
  \[92] ,
  \[16] ,
  \[93] ,
  \[17] ,
  \[94] ,
  MIS9174,
  \[18] ,
  \[95] ,
  \[19] ,
  \[96] ,
  \[97] ,
  \[98] ,
  \[20] ,
  MIS15328,
  \[21] ,
  \[22] ,
  \[23] ,
  MIS15339,
  \[24] ,
  \[25] ,
  MIS9255,
  \[26] ,
  \[27] ,
  \[28] ,
  \[29] ,
  MIS11546,
  MIS11547,
  MIS11548,
  MIS11549,
  MIS11560,
  MIS11562,
  MIS11565,
  MIS11550,
  MIS11556,
  MIS11581,
  MIS11582,
  MIS11583,
  MIS11584,
  MIS11585,
  MIS11586,
  MIS11587,
  MIS11588,
  MIS11589,
  \[30] ,
  MIS11578,
  \[31] ,
  MIS7401,
  \[32] ,
  MIS11590,
  MIS11591,
  MIS11592,
  MIS11593,
  MIS11594,
  \[33] ,
  \[34] ,
  \[35] ,
  \[36] ,
  \[37] ,
  MIS16602,
  MIS16604,
  MIS16606,
  MIS16609,
  MIS15650,
  \[38] ,
  \[39] ,
  MIS16620,
  MIS16623,
  MIS16625,
  MIS16627,
  MIS16629,
  MIS16611,
  MIS16613,
  MIS16615,
  MIS16618,
  MIS16646,
  MIS16631,
  MIS16633,
  MIS16665,
  MIS16657,
  \[40] ,
  MIS16670,
  MIS16673,
  MIS16675,
  \[41] ,
  \[42] ,
  MIS16690,
  \[43] ,
  \[44] ,
  \[45] ,
  \[46] ,
  \[47] ,
  MIS7564,
  \[48] ,
  \[49] ,
  MIS16541,
  MIS16544,
  MIS16546,
  MIS16548,
  MIS16565,
  MIS16569,
  MIS16553,
  MIS16555,
  MIS16581,
  MIS16583,
  MIS16585,
  MIS16588,
  \[50] ,
  MIS16572,
  MIS16577,
  MIS16579,
  \[51] ,
  \[52] ,
  MIS16591,
  MIS16593,
  MIS16596,
  MIS16598,
  \[53] ,
  MIS15062,
  MIS8641,
  MIS15065,
  \[54] ,
  MIS15843,
  \[55] ,
  MIS15847,
  MIS15848,
  MIS15080,
  MIS15081,
  MIS15083,
  \[56] ,
  MIS16023,
  MIS16027,
  \[57] ,
  \[58] ,
  MIS15854,
  MIS15855,
  \[59] ,
  MIS10125,
  MIS16864,
  MIS16866,
  MIS16858,
  MIS16883,
  MIS16885,
  MIS10130,
  MIS16887,
  MIS16889;
assign
  \[60]  = (MIS11590 & V1ZZZ4) | (MIS11589 & V1ZZZ3),
  MIS16871 = (~XZ163 & ~SLAD3) | (XZ163 & SLAD3),
  MIS16873 = (~SLAD2 & ~XZ162) | (SLAD2 & XZ162),
  MIS16879 = (XZFS & ~ICLR) | \[46] ,
  \[61]  = (MIS11590 & V1ZZZ5) | (MIS11589 & V1ZZZ4),
  V2ZZZ2_P = \[67] ,
  \[62]  = (MIS11590 & V1ZZZ6) | (MIS11589 & V1ZZZ5),
  MIS16891 = INZZZE | ~INYBB0,
  MIS16893 = ~VZZZE | ~VYBB0,
  MIS16895 = ~CBT2 | (CBT1 | CBT0),
  \[63]  = (MIS11590 & V1ZZZ7) | (MIS11589 & V1ZZZ6),
  QPR3_P = \[53] ,
  XZ323_P = \[92] ,
  \[64]  = (MIS11590 & VYBB1) | (MIS11589 & V1ZZZ7),
  P1ZZZ4_P = \[8] ,
  \[65]  = (MIS11592 & V2ZZZ1) | (MIS11591 & V2ZZZ0),
  I1ZZZ3_P = \[23] ,
  \[66]  = (MIS11592 & V2ZZZ2) | (MIS11591 & V2ZZZ1),
  TXWRD5_P = \[78] ,
  \[67]  = (MIS11592 & V2ZZZ3) | (MIS11591 & V2ZZZ2),
  MIS16701 = (MIS7401 & (TXWRD0 & MIS9255)) | (A & MIS16716),
  MIS16706 = (MIS16710 & (~QPR4 & (~QPR3 & MIS16690))) | ((MIS16712 & (RPTEN & RPTWIN)) | (~TXMESS_N & (MIS16701 & ~RPTWIN))),
  \[68]  = (MIS11592 & V2ZZZ4) | (MIS11591 & V2ZZZ3),
  MIS11154 = (MIS16690 & (~QPR4 & (~QPR3 & ~MIS9255))) | (TXWRD0 & MIS9255),
  STW_F = \[1] ,
  TXWRD13_P = \[86] ,
  \[69]  = (MIS11592 & V2ZZZ5) | (MIS11591 & V2ZZZ4),
  MIS16722 = (~MIS15650 & (~SLAD1 & ~SLAD0)) | ((MIS16724 & RPTWIN) | MIS15847),
  MIS16724 = ~RXZ1 | ~RXZ0,
  MIS16726 = (MIS11549 & TXWRD4) | ((MIS11548 & TXWRD3) | (V1ZZZ3 & VFIN)),
  MIS16728 = (MIS11549 & TXWRD5) | ((MIS11548 & TXWRD4) | (V1ZZZ4 & VFIN)),
  MIS16710 = (MIS7401 & (~MIS9255 & ~RPTWIN)) | ~\[0] ,
  MIS16712 = (~RXZ1 & (RXZ0 & ~ESRSUM)) | (RXZ1 & (~RXZ0 & ESRSUM)),
  MIS16716 = (~AXZ1 & (AXZ0 & ~MMERR)) | (AXZ1 & MIS16719),
  V1ZZZ4_P = \[61] ,
  MIS16719 = (~COMPPAR & AXZ0) | (~AXZ0 & ESRSUM),
  MIS16740 = (MIS11560 & MIS16742) | MIS15339,
  MIS16742 = ~XZ323 | ~XZ322,
  MIS16746 = (~MIS16767 & QPR3) | (~QPR3 & MIS16750),
  P2ZZZ1_P = \[13] ,
  MIS16748 = (~MIS16765 & ~TXMESS_N) | A,
  \[0]  = RPTWIN | ~TXMESS_N,
  MIS16730 = (MIS11560 & ~XZ322) | MIS15339,
  MIS16732 = (MIS11549 & TXWRD6) | ((MIS11548 & TXWRD5) | (V1ZZZ5 & VFIN)),
  MIS16734 = (MIS11549 & TXWRD14) | ((MIS11548 & TXWRD13) | (V2ZZZ5 & VFIN)),
  MIS16736 = (MIS11549 & TXWRD15) | ((MIS11548 & TXWRD14) | (V2ZZZ6 & VFIN)),
  I2ZZZ2_P = \[30] ,
  \[1]  = (MIS16790 & (MIS11547 & ~VFIN)) | RYZ,
  MIS16760 = (~TXMESS_N & (~QPR4 & (~QPR3 & (~B & (~MIS8768 & ~MIS15328))))) | (MIS16758 & B),
  MIS16762 = (~MIS9174 & ~C) | (MIS9174 & C),
  MIS16765 = ~MIS16746 | MIS8768,
  MIS16767 = ~B | QPR4,
  \[2]  = ~RYZ & MIS16706,
  MIS16750 = QPR4 | ~CBT2,
  MIS8768 = ~QPR2 | (QPR1 | ~QPR0),
  MIS16752 = MIS15847 | RPTWIN,
  MIS16754 = (MIS11560 & MIS7564) | \[89] ,
  MIS16758 = (~QPR3 & MIS15328) | (QPR4 | (MIS8768 | TXMESS_N)),
  \[3]  = (\[45]  & OFS2) | (XZFR1 & ~ICLR),
  MIS8027 = MIS7564 | (XZ163 | (XZ162 | (XZ161 | ~XZ160_N))),
  MIS16780 = (~QPR0 & SLAD1) | (QPR0 & SLAD0),
  MIS16786 = (\[46]  & XZFS) | (ENWIN & ~ICLR),
  MIS16788 = ~OFS1 | ~OFS2,
  TXWRD0_P = \[73] ,
  \[4]  = (MIS11588 & PYBB1) | (MIS11587 & P1ZZZ0),
  \[70]  = (MIS11592 & V2ZZZ6) | (MIS11591 & V2ZZZ5),
  A_P = \[47] ,
  MIS16778 = (SLAD3 & ~QPR0) | (SLAD2 & QPR0),
  \[5]  = (MIS11588 & PYBB2) | (MIS11587 & P1ZZZ1),
  \[71]  = (MIS11592 & V2ZZZ7) | (MIS11591 & V2ZZZ6),
  V2ZZZ1_P = \[66] ,
  \[6]  = (MIS11588 & PYBB3) | (MIS11587 & P1ZZZ2),
  \[72]  = (MIS11592 & VYBB1) | (MIS11591 & V2ZZZ7),
  MIS16790 = (MIS11556 & A) | STW_N,
  MIS16792 = ~MIS9255 | TXMESS_N,
  \[7]  = (MIS11588 & PYBB4) | (MIS11587 & P1ZZZ3),
  \[73]  = ~RYZ & MIS16591,
  TXWRD8_P = \[81] ,
  QPR4_P = \[54] ,
  XZ324_P = \[93] ,
  \[8]  = (MIS11588 & PYBB5) | (MIS11587 & P1ZZZ4),
  \[74]  = (MIS16606 & MIS11593) | (I1ZZZ1 & MIS11594),
  P1ZZZ3_P = \[7] ,
  \[9]  = (MIS11588 & PYBB6) | (MIS11587 & P1ZZZ5),
  \[75]  = (I1ZZZ2 & MIS11594) | (MIS16585 & MIS11593),
  I1ZZZ4_P = \[24] ,
  \[76]  = (MIS15080 & MIS16726) | ((P1ZZZ3 & MIS15081) | (I1ZZZ3 & MIS11594)),
  \[77]  = (MIS15080 & MIS16728) | ((P1ZZZ4 & MIS15081) | (I1ZZZ4 & MIS11594)),
  \[78]  = (MIS15080 & MIS16732) | ((P1ZZZ5 & MIS15081) | (I1ZZZ5 & MIS11594)),
  \[79]  = (MIS15080 & MIS16633) | ((P1ZZZ6 & MIS15081) | (I1ZZZ6 & MIS11594)),
  MIS12425 = MIS16673 | ~XZ320,
  V1ZZZ3_P = \[60] ,
  COMPPAR_P = \[38] ,
  XZFS_P = \[42] ,
  P2ZZZ4_P = \[16] ,
  I2ZZZ3_P = \[31] ,
  \[80]  = ~RYZ & MIS16618,
  XZ160_F = \[94] ,
  B_P = \[48] ,
  TXMESS_F = \[36] ,
  \[81]  = (MIS15080 & MIS16631) | ((P2ZZZ0 & MIS15081) | (I2ZZZ0 & MIS11594)),
  MIS9061 = (MIS16765 & ~A) | TXMESS_N,
  \[82]  = (MIS16627 & MIS11593) | (I2ZZZ1 & MIS11594),
  \[83]  = MIS16609 & ~RYZ,
  TXWRD7_P = \[80] ,
  MIS15964 = (MIS12425 & ~XZFS) | ((MIS16657 & SLAD0) | ((MIS16675 & MIS15650) | ((~PSYNC & MIS16673) | ((SLAD3 & MIS16665) | ((MIS16646 & SLAD1) | (SLAD2 & MIS16670)))))),
  \[84]  = ~RYZ & MIS16596,
  MIS9071 = (MIS11560 & MIS10125) | \[89] ,
  P1ZZZ6_P = \[10] ,
  V2ZZZ4_P = \[69] ,
  \[85]  = ~RYZ & MIS16623,
  I1ZZZ5_P = \[25] ,
  \[86]  = (MIS15080 & MIS16734) | ((I2ZZZ5 & MIS11594) | (P2ZZZ5 & MIS15081)),
  \[87]  = (MIS15080 & MIS16736) | ((I2ZZZ6 & MIS11594) | (P2ZZZ6 & MIS15081)),
  \[88]  = (MIS16583 & MIS11593) | (I2ZZZ7 & MIS11594),
  TXWRD15_P = \[88] ,
  \[89]  = MIS11560 & ~XZ320,
  V1ZZZ6_P = \[63] ,
  XZ161_P = \[95] ,
  RPTWIN_P = \[39] ,
  \[10]  = (MIS11588 & PYBB7) | (MIS11587 & P1ZZZ6),
  \[11]  = (MIS11588 & PYBB8) | (MIS11587 & P1ZZZ7),
  P2ZZZ3_P = \[15] ,
  \[12]  = (MIS11586 & PYBB1) | (MIS11585 & P2ZZZ0),
  AXZ0_P = \[55] ,
  I2ZZZ4_P = \[32] ,
  \[13]  = (MIS11586 & PYBB2) | (MIS11585 & P2ZZZ1),
  TXWRD2_P = \[75] ,
  \[90]  = (\[89]  & XZ321) | (MIS15083 & ~XZ321),
  C_P = \[49] ,
  \[14]  = (MIS11586 & PYBB3) | (MIS11585 & P2ZZZ2),
  \[91]  = (MIS15083 & (~XZ322 & XZ321)) | (MIS15339 & XZ322),
  \[15]  = (MIS11586 & PYBB4) | (MIS11585 & P2ZZZ3),
  \[92]  = (MIS11578 & (MIS15083 & ~XZ323)) | (MIS16730 & XZ323),
  \[16]  = (MIS11586 & PYBB5) | (MIS11585 & P2ZZZ4),
  \[93]  = (MIS11560 & (MIS11550 & ~XZ324)) | (MIS16740 & XZ324),
  \[17]  = (MIS11586 & PYBB6) | (MIS11585 & P2ZZZ5),
  \[94]  = (~MIS10125 & MIS15083) | (MIS16754 & XZ160_N),
  MIS9174 = (MIS16895 & ~QPR4) | (TXMESS_N | (QPR3 | MIS8768)),
  P1ZZZ5_P = \[9] ,
  V2ZZZ3_P = \[68] ,
  \[18]  = (MIS11586 & PYBB7) | (MIS11585 & P2ZZZ6),
  \[95]  = (MIS15083 & (~MIS10125 & ~XZ161)) | (MIS9071 & XZ161),
  I1ZZZ6_P = \[26] ,
  \[19]  = (MIS11586 & PYBB8) | (MIS11585 & P2ZZZ7),
  \[96]  = (MIS11560 & (~XZ162 & MIS15848)) | (XZ162 & MIS16588),
  \[97]  = (MIS11560 & (~XZ163 & (XZ162 & MIS15848))) | (MIS16602 & XZ163),
  FSESR_P = \[3] ,
  \[98]  = MIS16788 & (MIS16786 & PSRW),
  V1ZZZ5_P = \[62] ,
  XZ162_P = \[96] ,
  TXWRD10_P = \[83] ,
  \[20]  = (MIS11582 & INYBB1) | (MIS11581 & I1ZZZ0),
  MIS15328 = (~CBT1 & ~CBT0) | ~CBT2,
  \[21]  = (MIS11582 & INYBB2) | (MIS11581 & I1ZZZ1),
  P1ZZZ0_P = \[4] ,
  OFS1_P = \[46] ,
  P2ZZZ6_P = \[18] ,
  \[22]  = (MIS11582 & INYBB3) | (MIS11581 & I1ZZZ2),
  AXZ1_P = \[56] ,
  I2ZZZ5_P = \[33] ,
  \[23]  = (MIS11582 & INYBB4) | (MIS11581 & I1ZZZ3),
  TXWRD1_P = \[74] ,
  MIS15339 = (MIS11560 & ~XZ321) | \[89] ,
  \[24]  = (MIS11582 & INYBB5) | (MIS11581 & I1ZZZ4),
  \[25]  = (MIS11582 & INYBB6) | (MIS11581 & I1ZZZ5),
  MIS9255 = C | B,
  I1ZZZ7_P = \[27] ,
  \[26]  = (MIS11582 & INYBB7) | (MIS11581 & I1ZZZ6),
  TXWRD9_P = \[82] ,
  ENWIN_P = \[98] ,
  \[27]  = (MIS11582 & INYBB8) | (MIS11581 & I1ZZZ7),
  V1ZZZ0_P = \[57] ,
  V2ZZZ6_P = \[71] ,
  \[28]  = (MIS11584 & INYBB1) | (MIS11583 & I2ZZZ0),
  \[29]  = (MIS11584 & INYBB2) | (MIS11583 & I2ZZZ1),
  MIS11546 = ~INFIN & PFIN,
  MIS11547 = ~INFIN & ~PFIN,
  MIS11548 = MIS16792 & ~VFIN,
  MIS11549 = ~MIS16792 & ~VFIN,
  MIS11560 = ~ICLR & ~PSYNC,
  MIS11562 = ~PFIN & VFIN,
  MIS11565 = MIS11547 & (~VFIN & TXMESS_N),
  XZ163_P = \[97] ,
  MIS11550 = MIS11578 & (XZ323 & XZ320),
  MIS11556 = AXZ1 & (AXZ0 & ~TXMESS_N),
  MIS11581 = ~RYZ & MIS16891,
  MIS11582 = ~MIS16891 & ~RYZ,
  MIS11583 = ~RYZ & MIS16887,
  MIS11584 = ~MIS16887 & ~RYZ,
  MIS11585 = ~RYZ & MIS16885,
  MIS11586 = ~MIS16885 & ~RYZ,
  MIS11587 = ~RYZ & MIS16883,
  MIS11588 = ~MIS16883 & ~RYZ,
  MIS11589 = ~RYZ & MIS16889,
  \[30]  = (MIS11584 & INYBB3) | (MIS11583 & I2ZZZ2),
  MIS11578 = XZ322 & XZ321,
  \[31]  = (MIS11584 & INYBB4) | (MIS11583 & I2ZZZ3),
  MIS7401 = (~AXZ1 & ~AXZ0) | ~A,
  OFS2_P = \[45] ,
  P2ZZZ5_P = \[17] ,
  \[32]  = (MIS11584 & INYBB5) | (MIS11583 & I2ZZZ4),
  MIS11590 = ~MIS16889 & ~RYZ,
  MIS11591 = ~RYZ & MIS16893,
  I1ZZZ0_P = \[20] ,
  MIS11592 = ~MIS16893 & ~RYZ,
  MIS11593 = ~RYZ & ~INFIN,
  MIS11594 = ~RYZ & INFIN,
  I2ZZZ6_P = \[34] ,
  \[33]  = (MIS11584 & INYBB6) | (MIS11583 & I2ZZZ5),
  QPR0_P = \[50] ,
  XZ320_P = \[89] ,
  \[34]  = (MIS11584 & INYBB7) | (MIS11583 & I2ZZZ6),
  P1ZZZ7_P = \[11] ,
  \[35]  = (MIS11584 & INYBB8) | (MIS11583 & I2ZZZ7),
  \[36]  = MIS11565 | RYZ,
  TXWRD4_P = \[77] ,
  RXZ0_P = \[43] ,
  \[37]  = (MIS11556 & A) | ICLR,
  MIS16602 = (MIS16604 & MIS11560) | MIS9071,
  MIS16604 = ~XZ161 | ~XZ162,
  MIS16606 = (MIS11562 & V1ZZZ1) | ((MIS15065 & TXWRD2) | ((MIS15062 & TXWRD1) | (P1ZZZ1 & PFIN))),
  MIS16609 = (I2ZZZ2 & INFIN) | ((MIS11547 & MIS16611) | (MIS11546 & P2ZZZ2)),
  MIS15650 = ~XZFS | (~PSYNC | (SLAD3 | SLAD2)),
  V2ZZZ5_P = \[70] ,
  \[38]  = ~RYZ & MIS16569,
  \[39]  = ~RYZ & MIS16722,
  MIS16620 = (MIS11549 & TXWRD8) | ((MIS11548 & TXWRD7) | (V1ZZZ7 & VFIN)),
  MIS16623 = (I2ZZZ4 & INFIN) | ((MIS16625 & MIS11547) | (MIS11546 & P2ZZZ4)),
  MIS16625 = (MIS11549 & TXWRD13) | ((MIS11548 & TXWRD12) | (V2ZZZ4 & VFIN)),
  SBUFF = \[0] ,
  MIS16627 = (MIS11562 & V2ZZZ1) | ((MIS15065 & TXWRD10) | ((MIS15062 & TXWRD9) | (P2ZZZ1 & PFIN))),
  MIS16629 = MIS11565 | ~QPR0,
  MIS16611 = (MIS11549 & TXWRD11) | ((MIS11548 & TXWRD10) | (V2ZZZ2 & VFIN)),
  MIS16613 = (MIS11560 & ~XZFR0) | MIS10130,
  MIS16615 = (~MIS9061 & ~AXZ0) | (MIS9061 & AXZ0),
  V1ZZZ7_P = \[64] ,
  MIS16618 = (P1ZZZ7 & MIS11546) | ((I1ZZZ7 & INFIN) | (MIS16620 & MIS11547)),
  MIS16646 = ~ENWIN | (~XZ161 | (MIS12425 | MIS16023)),
  P2ZZZ0_P = \[12] ,
  MIS16631 = (MIS11549 & TXWRD9) | ((MIS11548 & TXWRD8) | (V2ZZZ0 & VFIN)),
  MIS16633 = (MIS11549 & TXWRD7) | ((MIS11548 & TXWRD6) | (V1ZZZ6 & VFIN)),
  MIS16665 = ~XZ320 | (MIS15855 | ~XZ163),
  MIS16657 = MIS12425 | (MIS16027 | MIS10125),
  TXWRD12_P = \[85] ,
  I2ZZZ7_P = \[35] ,
  \[40]  = (MIS15083 & (~MIS8027 & ~XZFR0)) | (MIS10130 & XZFR0),
  MIS16670 = ~XZ320 | (MIS15854 | ~XZ162),
  MIS16673 = MIS15855 | MIS15854,
  MIS16675 = MIS16027 | MIS16023,
  \[41]  = (~MIS8027 & (MIS15083 & (~XZFR1 & XZFR0))) | (MIS16613 & XZFR1),
  P1ZZZ2_P = \[6] ,
  V2ZZZ0_P = \[65] ,
  \[42]  = MIS16788 & (MIS16879 & PSRW),
  MIS16690 = (MIS16780 & (QPR2 & ~QPR1)) | (MIS16778 & (~QPR2 & QPR1)),
  I1ZZZ1_P = \[21] ,
  \[43]  = (MIS16544 & (RXZ0 & ~RPTWIN)) | (MIS8641 & ~RXZ0),
  QPR1_P = \[51] ,
  XZ321_P = \[90] ,
  \[44]  = (MIS8641 & (~RXZ1 & RXZ0)) | (MIS16541 & RXZ1),
  \[45]  = OFS1 & ~ICLR,
  \[46]  = ~ICLR & PSYNC,
  TXWRD3_P = \[76] ,
  RXZ1_P = \[44] ,
  \[47]  = ~RYZ & MIS16748,
  V1ZZZ2_P = \[59] ,
  MIS7564 = ~MIS11578 | (~XZ324 | ~XZ323),
  XZFR0_P = \[40] ,
  TD_P = \[2] ,
  \[48]  = ~RYZ & MIS16760,
  \[49]  = ~RYZ & MIS16762,
  MIS16541 = (~ICLR & ~RXZ0) | (MIS16544 & ~RPTWIN),
  MIS16544 = (MIS15964 & ~ICLR) | \[89] ,
  MIS16546 = MIS16548 | ~QPR3,
  MIS16548 = MIS16581 | ~QPR2,
  I2ZZZ0_P = \[28] ,
  MIS16565 = (~COMPPAR & (~TXMESS_N & MIS16577)) | ((COMPPAR & MIS16579) | MIS11556),
  MIS16569 = (~COMPPAR & (~TXMESS_N & (MIS7401 & MIS11154))) | ((COMPPAR & MIS16572) | (A & MIS16565)),
  MIS16553 = (~AXZ1 & (AXZ0 & ~MIS9061)) | (MIS16555 & AXZ1),
  MIS16555 = ~AXZ0 | MIS9061,
  P2ZZZ7_P = \[19] ,
  TXWRD11_P = \[84] ,
  MIS16581 = MIS16629 | ~QPR1,
  MIS16583 = (MIS11562 & V2ZZZ7) | ((MIS15062 & TXWRD15) | (P2ZZZ7 & PFIN)),
  MIS16585 = (MIS11562 & V1ZZZ2) | ((MIS15065 & TXWRD3) | ((MIS15062 & TXWRD2) | (P1ZZZ2 & PFIN))),
  MIS16588 = (MIS11560 & ~XZ161) | MIS9071,
  \[50]  = (MIS11565 & (QPR0 & ~RYZ)) | (~\[36]  & ~QPR0),
  MIS16572 = (MIS7401 & ~MIS11154) | TXMESS_N,
  MIS16577 = (AXZ1 & ESRSUM) | (AXZ0 & ~MMERR),
  MIS16579 = (AXZ1 & ~ESRSUM) | (AXZ0 & MMERR),
  \[51]  = (~RYZ & (MIS16629 & QPR1)) | (~\[36]  & (~QPR1 & QPR0)),
  P1ZZZ1_P = \[5] ,
  \[52]  = (~RYZ & (MIS16581 & QPR2)) | (MIS15843 & ~QPR2),
  MIS16591 = (P1ZZZ0 & MIS11546) | ((MIS16593 & MIS11547) | (I1ZZZ0 & INFIN)),
  MIS16593 = (MIS11549 & TXWRD1) | ((MIS11548 & TXWRD0) | (V1ZZZ0 & VFIN)),
  I1ZZZ2_P = \[22] ,
  MIS16596 = (I2ZZZ3 & INFIN) | ((MIS16598 & MIS11547) | (MIS11546 & P2ZZZ3)),
  MIS16598 = (MIS11549 & TXWRD12) | ((MIS11548 & TXWRD11) | (V2ZZZ3 & VFIN)),
  RYZ_P = \[37] ,
  \[53]  = (~RYZ & (MIS16548 & QPR3)) | (MIS15843 & (~QPR3 & QPR2)),
  QPR2_P = \[52] ,
  XZ322_P = \[91] ,
  MIS15062 = MIS11548 & ~PFIN,
  MIS8641 = (~SLAD3 & (~SLAD2 & (~SLAD1 & (~SLAD0 & (XZFS & \[46] ))))) | (~ICLR & MIS16752),
  MIS15065 = MIS11549 & ~PFIN,
  \[54]  = (MIS15843 & (~QPR4 & (QPR3 & QPR2))) | (~RYZ & (QPR4 & MIS16546)),
  V2ZZZ7_P = \[72] ,
  MIS15843 = ~\[36]  & (QPR0 & QPR1),
  \[55]  = ~RYZ & MIS16615,
  MIS15847 = MIS16866 & (MIS16864 & (MIS16858 & (MIS11550 & (ENWIN & XZ324)))),
  MIS15848 = ~MIS10125 & (XZ161 & XZ320),
  MIS15080 = MIS11593 & ~PFIN,
  MIS15081 = MIS11593 & PFIN,
  MIS15083 = MIS11560 & XZ320,
  \[56]  = ~RYZ & MIS16553,
  MIS16023 = (~XZ160_N & ~SLAD0) | MIS7564,
  TXWRD6_P = \[79] ,
  MIS16027 = (XZ161 & ~SLAD1) | ~ENWIN,
  \[57]  = (MIS11590 & V1ZZZ1) | (MIS11589 & V1ZZZ0),
  V1ZZZ1_P = \[58] ,
  XZFR1_P = \[41] ,
  \[58]  = (MIS11590 & V1ZZZ2) | (MIS11589 & V1ZZZ1),
  MIS15854 = XZ163 & ~SLAD3,
  MIS15855 = XZ162 & ~SLAD2,
  TXWRD14_P = \[87] ,
  \[59]  = (MIS11590 & V1ZZZ3) | (MIS11589 & V1ZZZ2),
  P2ZZZ2_P = \[14] ,
  I2ZZZ1_P = \[29] ,
  MIS10125 = MIS7564 | XZ160_N,
  MIS16864 = (~SLAD1 & ~XZ161) | (SLAD1 & XZ161),
  MIS16866 = (~SLAD0 & XZ160_N) | (SLAD0 & ~XZ160_N),
  MIS16858 = MIS16873 & MIS16871,
  MIS16883 = PZZZE | ~PYBB0,
  MIS16885 = ~PZZZE | ~PYBB0,
  MIS10130 = (MIS11560 & MIS8027) | \[89] ,
  MIS16887 = ~INZZZE | ~INYBB0,
  MIS16889 = VZZZE | ~VYBB0;
endmodule

