// C6288
module foobar(g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x, y, z, a0, b0, c0, d0, e0, f0);
input a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x, y, z, a0, b0, c0, d0, e0, f0;
output g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1;
and(g0, a, q);
not(t_0, b17);
not(t_1, c17);
and(h0, t_0, t_1);
not(t_2, f22);
not(t_3, i22);
and(i0, t_2, t_3);
not(t_4, l27);
not(t_5, q27);
and(j0, t_4, t_5);
not(t_6, s32);
not(t_7, z32);
and(k0, t_6, t_7);
not(t_8, a38);
not(t_9, j38);
and(l0, t_8, t_9);
not(t_10, l43);
not(t_11, w43);
and(m0, t_10, t_11);
not(t_12, y48);
not(t_13, l49);
and(n0, t_12, t_13);
not(t_14, n54);
not(t_15, c55);
and(o0, t_14, t_15);
not(t_16, g60);
not(t_17, u60);
and(p0, t_16, t_17);
not(t_18, a66);
not(t_19, n66);
and(q0, t_18, t_19);
not(t_20, x71);
not(t_21, j72);
and(r0, t_20, t_21);
not(t_22, x77);
not(t_23, h78);
and(s0, t_22, t_23);
not(t_24, x83);
not(t_25, h84);
and(t0, t_24, t_25);
not(t_26, a89);
not(t_27, g89);
and(u0, t_26, t_27);
not(t_28, s91);
not(t_29, u91);
and(v0, t_28, t_29);
not(t_30, f92);
not(t_31, g92);
and(w0, t_30, t_31);
not(t_32, j92);
not(t_33, k92);
and(x0, t_32, t_33);
not(t_34, n92);
not(t_35, o92);
and(y0, t_34, t_35);
not(t_36, r92);
not(t_37, s92);
and(z0, t_36, t_37);
not(t_38, v92);
not(t_39, w92);
and(a1, t_38, t_39);
not(t_40, z92);
not(t_41, a93);
and(b1, t_40, t_41);
not(t_42, d93);
not(t_43, e93);
and(c1, t_42, t_43);
not(t_44, h93);
not(t_45, i93);
and(d1, t_44, t_45);
not(t_46, l93);
not(t_47, m93);
and(e1, t_46, t_47);
not(t_48, p93);
not(t_49, q93);
and(f1, t_48, t_49);
not(t_50, t93);
not(t_51, u93);
and(g1, t_50, t_51);
not(t_52, x93);
not(t_53, y93);
and(h1, t_52, t_53);
not(t_54, b94);
not(t_55, c94);
and(i1, t_54, t_55);
not(t_56, f94);
not(t_57, g94);
and(j1, t_56, t_57);
not(t_58, d82);
not(t_59, h94);
and(k1, t_58, t_59);
not(t_60, i94);
not(t_61, j94);
and(l1, t_60, t_61);
and(s2, p, f0);
and(t2, p, e0);
and(u2, p, d0);
and(v2, p, c0);
and(w2, p, b0);
and(x2, p, a0);
and(y2, p, z);
and(z2, p, y);
and(a3, p, x);
and(b3, p, w);
and(c3, p, v);
and(d3, p, u);
and(e3, p, t);
and(f3, p, s);
and(g3, p, r);
and(h3, p, q);
and(i3, o, f0);
and(j3, o, e0);
and(k3, o, d0);
and(l3, o, c0);
and(m3, o, b0);
and(n3, o, a0);
and(o3, o, z);
and(p3, o, y);
and(q3, o, x);
and(r3, o, w);
and(s3, o, v);
and(t3, o, u);
and(u3, o, t);
and(v3, o, s);
and(w3, o, r);
and(x3, o, q);
and(y3, n, f0);
and(z3, n, e0);
and(a4, n, d0);
and(b4, n, c0);
and(c4, n, b0);
and(d4, n, a0);
and(e4, n, z);
and(f4, n, y);
and(g4, n, x);
and(h4, n, w);
and(i4, n, v);
and(j4, n, u);
and(k4, n, t);
and(l4, n, s);
and(m4, n, r);
and(n4, n, q);
and(o4, m, f0);
and(p4, m, e0);
and(q4, m, d0);
and(r4, m, c0);
and(s4, m, b0);
and(t4, m, a0);
and(u4, m, z);
and(v4, m, y);
and(w4, m, x);
and(x4, m, w);
and(y4, m, v);
and(z4, m, u);
and(a5, m, t);
and(b5, m, s);
and(c5, m, r);
and(d5, m, q);
and(e5, l, f0);
and(f5, l, e0);
and(g5, l, d0);
and(h5, l, c0);
and(i5, l, b0);
and(j5, l, a0);
and(k5, l, z);
and(l5, l, y);
and(m5, l, x);
and(n5, l, w);
and(o5, l, v);
and(p5, l, u);
and(q5, l, t);
and(r5, l, s);
and(s5, l, r);
and(t5, l, q);
and(u5, k, f0);
and(v5, k, e0);
and(w5, k, d0);
and(x5, k, c0);
and(y5, k, b0);
and(z5, k, a0);
and(a6, k, z);
and(b6, k, y);
and(c6, k, x);
and(d6, k, w);
and(e6, k, v);
and(f6, k, u);
and(g6, k, t);
and(h6, k, s);
and(i6, k, r);
and(j6, k, q);
and(k6, j, f0);
and(l6, j, e0);
and(m6, j, d0);
and(n6, j, c0);
and(o6, j, b0);
and(p6, j, a0);
and(q6, j, z);
and(r6, j, y);
and(s6, j, x);
and(t6, j, w);
and(u6, j, v);
and(v6, j, u);
and(w6, j, t);
and(x6, j, s);
and(y6, j, r);
and(z6, j, q);
and(a7, i, f0);
and(b7, i, e0);
and(c7, i, d0);
and(d7, i, c0);
and(e7, i, b0);
and(f7, i, a0);
and(g7, i, z);
and(h7, i, y);
and(i7, i, x);
and(j7, i, w);
and(k7, i, v);
and(l7, i, u);
and(m7, i, t);
and(n7, i, s);
and(o7, i, r);
and(p7, i, q);
and(q7, h, f0);
and(r7, h, e0);
and(s7, h, d0);
and(t7, h, c0);
and(u7, h, b0);
and(v7, h, a0);
and(w7, h, z);
and(x7, h, y);
and(y7, h, x);
and(z7, h, w);
and(a8, h, v);
and(b8, h, u);
and(c8, h, t);
and(d8, h, s);
and(e8, h, r);
and(f8, h, q);
and(g8, g, f0);
and(h8, g, e0);
and(i8, g, d0);
and(j8, g, c0);
and(k8, g, b0);
and(l8, g, a0);
and(m8, g, z);
and(n8, g, y);
and(o8, g, x);
and(p8, g, w);
and(q8, g, v);
and(r8, g, u);
and(s8, g, t);
and(t8, g, s);
and(u8, g, r);
and(v8, g, q);
and(w8, f, f0);
and(x8, f, e0);
and(y8, f, d0);
and(z8, f, c0);
and(a9, f, b0);
and(b9, f, a0);
and(c9, f, z);
and(d9, f, y);
and(e9, f, x);
and(f9, f, w);
and(g9, f, v);
and(h9, f, u);
and(i9, f, t);
and(j9, f, s);
and(k9, f, r);
and(l9, f, q);
and(m9, e, f0);
and(n9, e, e0);
and(o9, e, d0);
and(p9, e, c0);
and(q9, e, b0);
and(r9, e, a0);
and(s9, e, z);
and(t9, e, y);
and(u9, e, x);
and(v9, e, w);
and(w9, e, v);
and(x9, e, u);
and(y9, e, t);
and(z9, e, s);
and(a10, e, r);
and(b10, e, q);
and(c10, d, f0);
and(d10, d, e0);
and(e10, d, d0);
and(f10, d, c0);
and(g10, d, b0);
and(h10, d, a0);
and(i10, d, z);
and(j10, d, y);
and(k10, d, x);
and(l10, d, w);
and(m10, d, v);
and(n10, d, u);
and(o10, d, t);
and(p10, d, s);
and(q10, d, r);
and(r10, d, q);
and(s10, c, f0);
and(t10, c, e0);
and(u10, c, d0);
and(v10, c, c0);
and(w10, c, b0);
and(x10, c, a0);
and(y10, c, z);
and(z10, c, y);
and(a11, c, x);
and(b11, c, w);
and(c11, c, v);
and(d11, c, u);
and(e11, c, t);
and(f11, c, s);
and(g11, c, r);
and(h11, c, q);
and(i11, b, f0);
and(j11, b, e0);
and(k11, b, d0);
and(l11, b, c0);
and(m11, b, b0);
and(n11, b, a0);
and(o11, b, z);
and(p11, b, y);
and(q11, b, x);
and(r11, b, w);
and(s11, b, v);
and(t11, b, u);
and(u11, b, t);
and(v11, b, s);
and(w11, b, r);
and(x11, b, q);
and(y11, a, f0);
and(z11, a, e0);
and(a12, a, d0);
and(b12, a, c0);
and(c12, a, b0);
and(d12, a, a0);
and(e12, a, z);
and(f12, a, y);
and(g12, a, x);
and(h12, a, w);
and(i12, a, v);
and(j12, a, u);
and(k12, a, t);
and(l12, a, s);
and(m12, a, r);
not(n12, h3);
not(o12, x3);
not(p12, n4);
not(q12, d5);
not(r12, t5);
not(s12, j6);
not(t12, z6);
not(u12, p7);
not(v12, f8);
not(w12, v8);
not(x12, l9);
not(y12, b10);
not(z12, r10);
not(a13, h11);
not(b13, x11);
not(c13, n12);
not(t_62, h3);
not(t_63, n12);
and(d13, t_62, t_63);
not(e13, o12);
not(t_64, x3);
not(t_65, o12);
and(f13, t_64, t_65);
not(g13, p12);
not(t_66, n4);
not(t_67, p12);
and(h13, t_66, t_67);
not(i13, q12);
not(t_68, d5);
not(t_69, q12);
and(j13, t_68, t_69);
not(k13, r12);
not(t_70, t5);
not(t_71, r12);
and(l13, t_70, t_71);
not(m13, s12);
not(t_72, j6);
not(t_73, s12);
and(n13, t_72, t_73);
not(o13, t12);
not(t_74, z6);
not(t_75, t12);
and(p13, t_74, t_75);
not(q13, u12);
not(t_76, p7);
not(t_77, u12);
and(r13, t_76, t_77);
not(s13, v12);
not(t_78, f8);
not(t_79, v12);
and(t13, t_78, t_79);
not(u13, w12);
not(t_80, v8);
not(t_81, w12);
and(v13, t_80, t_81);
not(w13, x12);
not(t_82, l9);
not(t_83, x12);
and(x13, t_82, t_83);
not(y13, y12);
not(t_84, b10);
not(t_85, y12);
and(z13, t_84, t_85);
not(a14, z12);
not(t_86, r10);
not(t_87, z12);
and(b14, t_86, t_87);
not(c14, a13);
not(t_88, h11);
not(t_89, a13);
and(d14, t_88, t_89);
not(e14, b13);
not(t_90, x11);
not(t_91, b13);
and(f14, t_90, t_91);
not(t_92, d13);
not(t_93, c13);
and(g14, t_92, t_93);
not(t_94, f13);
not(t_95, e13);
and(h14, t_94, t_95);
not(t_96, h13);
not(t_97, g13);
and(i14, t_96, t_97);
not(t_98, j13);
not(t_99, i13);
and(j14, t_98, t_99);
not(t_100, l13);
not(t_101, k13);
and(k14, t_100, t_101);
not(t_102, n13);
not(t_103, m13);
and(l14, t_102, t_103);
not(t_104, p13);
not(t_105, o13);
and(m14, t_104, t_105);
not(t_106, r13);
not(t_107, q13);
and(n14, t_106, t_107);
not(t_108, t13);
not(t_109, s13);
and(o14, t_108, t_109);
not(t_110, v13);
not(t_111, u13);
and(p14, t_110, t_111);
not(t_112, x13);
not(t_113, w13);
and(q14, t_112, t_113);
not(t_114, z13);
not(t_115, y13);
and(r14, t_114, t_115);
not(t_116, b14);
not(t_117, a14);
and(s14, t_116, t_117);
not(t_118, d14);
not(t_119, c14);
and(t14, t_118, t_119);
not(t_120, f14);
not(t_121, e14);
and(u14, t_120, t_121);
not(t_122, g14);
not(t_123, w3);
and(v14, t_122, t_123);
not(t_124, h14);
not(t_125, m4);
and(w14, t_124, t_125);
not(t_126, i14);
not(t_127, c5);
and(x14, t_126, t_127);
not(t_128, j14);
not(t_129, s5);
and(y14, t_128, t_129);
not(t_130, k14);
not(t_131, i6);
and(z14, t_130, t_131);
not(t_132, l14);
not(t_133, y6);
and(a15, t_132, t_133);
not(t_134, m14);
not(t_135, o7);
and(b15, t_134, t_135);
not(t_136, n14);
not(t_137, e8);
and(c15, t_136, t_137);
not(t_138, o14);
not(t_139, u8);
and(d15, t_138, t_139);
not(t_140, p14);
not(t_141, k9);
and(e15, t_140, t_141);
not(t_142, q14);
not(t_143, a10);
and(f15, t_142, t_143);
not(t_144, r14);
not(t_145, q10);
and(g15, t_144, t_145);
not(t_146, s14);
not(t_147, g11);
and(h15, t_146, t_147);
not(t_148, t14);
not(t_149, w11);
and(i15, t_148, t_149);
not(t_150, u14);
not(t_151, m12);
and(j15, t_150, t_151);
not(t_152, n12);
not(t_153, v14);
and(k15, t_152, t_153);
not(t_154, g14);
not(t_155, v14);
and(l15, t_154, t_155);
not(t_156, v14);
not(t_157, w3);
and(m15, t_156, t_157);
not(t_158, o12);
not(t_159, w14);
and(n15, t_158, t_159);
not(t_160, h14);
not(t_161, w14);
and(o15, t_160, t_161);
not(t_162, w14);
not(t_163, m4);
and(p15, t_162, t_163);
not(t_164, p12);
not(t_165, x14);
and(q15, t_164, t_165);
not(t_166, i14);
not(t_167, x14);
and(r15, t_166, t_167);
not(t_168, x14);
not(t_169, c5);
and(s15, t_168, t_169);
not(t_170, q12);
not(t_171, y14);
and(t15, t_170, t_171);
not(t_172, j14);
not(t_173, y14);
and(u15, t_172, t_173);
not(t_174, y14);
not(t_175, s5);
and(v15, t_174, t_175);
not(t_176, r12);
not(t_177, z14);
and(w15, t_176, t_177);
not(t_178, k14);
not(t_179, z14);
and(x15, t_178, t_179);
not(t_180, z14);
not(t_181, i6);
and(y15, t_180, t_181);
not(t_182, s12);
not(t_183, a15);
and(z15, t_182, t_183);
not(t_184, l14);
not(t_185, a15);
and(a16, t_184, t_185);
not(t_186, a15);
not(t_187, y6);
and(b16, t_186, t_187);
not(t_188, t12);
not(t_189, b15);
and(c16, t_188, t_189);
not(t_190, m14);
not(t_191, b15);
and(d16, t_190, t_191);
not(t_192, b15);
not(t_193, o7);
and(e16, t_192, t_193);
not(t_194, u12);
not(t_195, c15);
and(f16, t_194, t_195);
not(t_196, n14);
not(t_197, c15);
and(g16, t_196, t_197);
not(t_198, c15);
not(t_199, e8);
and(h16, t_198, t_199);
not(t_200, v12);
not(t_201, d15);
and(i16, t_200, t_201);
not(t_202, o14);
not(t_203, d15);
and(j16, t_202, t_203);
not(t_204, d15);
not(t_205, u8);
and(k16, t_204, t_205);
not(t_206, w12);
not(t_207, e15);
and(l16, t_206, t_207);
not(t_208, p14);
not(t_209, e15);
and(m16, t_208, t_209);
not(t_210, e15);
not(t_211, k9);
and(n16, t_210, t_211);
not(t_212, x12);
not(t_213, f15);
and(o16, t_212, t_213);
not(t_214, q14);
not(t_215, f15);
and(p16, t_214, t_215);
not(t_216, f15);
not(t_217, a10);
and(q16, t_216, t_217);
not(t_218, y12);
not(t_219, g15);
and(r16, t_218, t_219);
not(t_220, r14);
not(t_221, g15);
and(s16, t_220, t_221);
not(t_222, g15);
not(t_223, q10);
and(t16, t_222, t_223);
not(t_224, z12);
not(t_225, h15);
and(u16, t_224, t_225);
not(t_226, s14);
not(t_227, h15);
and(v16, t_226, t_227);
not(t_228, h15);
not(t_229, g11);
and(w16, t_228, t_229);
not(t_230, a13);
not(t_231, i15);
and(x16, t_230, t_231);
not(t_232, t14);
not(t_233, i15);
and(y16, t_232, t_233);
not(t_234, i15);
not(t_235, w11);
and(z16, t_234, t_235);
not(t_236, b13);
not(t_237, j15);
and(a17, t_236, t_237);
not(t_238, u14);
not(t_239, j15);
and(b17, t_238, t_239);
not(t_240, j15);
not(t_241, m12);
and(c17, t_240, t_241);
not(t_242, g3);
not(t_243, k15);
and(d17, t_242, t_243);
not(t_244, l15);
not(t_245, m15);
and(e17, t_244, t_245);
not(t_246, o15);
not(t_247, p15);
and(f17, t_246, t_247);
not(t_248, r15);
not(t_249, s15);
and(g17, t_248, t_249);
not(t_250, u15);
not(t_251, v15);
and(h17, t_250, t_251);
not(t_252, x15);
not(t_253, y15);
and(i17, t_252, t_253);
not(t_254, a16);
not(t_255, b16);
and(j17, t_254, t_255);
not(t_256, d16);
not(t_257, e16);
and(k17, t_256, t_257);
not(t_258, g16);
not(t_259, h16);
and(l17, t_258, t_259);
not(t_260, j16);
not(t_261, k16);
and(m17, t_260, t_261);
not(t_262, m16);
not(t_263, n16);
and(n17, t_262, t_263);
not(t_264, p16);
not(t_265, q16);
and(o17, t_264, t_265);
not(t_266, s16);
not(t_267, t16);
and(p17, t_266, t_267);
not(t_268, v16);
not(t_269, w16);
and(q17, t_268, t_269);
not(t_270, y16);
not(t_271, z16);
and(r17, t_270, t_271);
not(t_272, g3);
not(t_273, d17);
and(s17, t_272, t_273);
not(t_274, d17);
not(t_275, k15);
and(t17, t_274, t_275);
not(t_276, e17);
not(t_277, n15);
and(u17, t_276, t_277);
not(t_278, f17);
not(t_279, q15);
and(v17, t_278, t_279);
not(t_280, g17);
not(t_281, t15);
and(w17, t_280, t_281);
not(t_282, h17);
not(t_283, w15);
and(x17, t_282, t_283);
not(t_284, i17);
not(t_285, z15);
and(y17, t_284, t_285);
not(t_286, j17);
not(t_287, c16);
and(z17, t_286, t_287);
not(t_288, k17);
not(t_289, f16);
and(a18, t_288, t_289);
not(t_290, l17);
not(t_291, i16);
and(b18, t_290, t_291);
not(t_292, m17);
not(t_293, l16);
and(c18, t_292, t_293);
not(t_294, n17);
not(t_295, o16);
and(d18, t_294, t_295);
not(t_296, o17);
not(t_297, r16);
and(e18, t_296, t_297);
not(t_298, p17);
not(t_299, u16);
and(f18, t_298, t_299);
not(t_300, q17);
not(t_301, x16);
and(g18, t_300, t_301);
not(t_302, r17);
not(t_303, a17);
and(h18, t_302, t_303);
not(t_304, s17);
not(t_305, t17);
and(i18, t_304, t_305);
not(t_306, e17);
not(t_307, u17);
and(j18, t_306, t_307);
not(t_308, u17);
not(t_309, n15);
and(k18, t_308, t_309);
not(t_310, f17);
not(t_311, v17);
and(l18, t_310, t_311);
not(t_312, v17);
not(t_313, q15);
and(m18, t_312, t_313);
not(t_314, g17);
not(t_315, w17);
and(n18, t_314, t_315);
not(t_316, w17);
not(t_317, t15);
and(o18, t_316, t_317);
not(t_318, h17);
not(t_319, x17);
and(p18, t_318, t_319);
not(t_320, x17);
not(t_321, w15);
and(q18, t_320, t_321);
not(t_322, i17);
not(t_323, y17);
and(r18, t_322, t_323);
not(t_324, y17);
not(t_325, z15);
and(s18, t_324, t_325);
not(t_326, j17);
not(t_327, z17);
and(t18, t_326, t_327);
not(t_328, z17);
not(t_329, c16);
and(u18, t_328, t_329);
not(t_330, k17);
not(t_331, a18);
and(v18, t_330, t_331);
not(t_332, a18);
not(t_333, f16);
and(w18, t_332, t_333);
not(t_334, l17);
not(t_335, b18);
and(x18, t_334, t_335);
not(t_336, b18);
not(t_337, i16);
and(y18, t_336, t_337);
not(t_338, m17);
not(t_339, c18);
and(z18, t_338, t_339);
not(t_340, c18);
not(t_341, l16);
and(a19, t_340, t_341);
not(t_342, n17);
not(t_343, d18);
and(b19, t_342, t_343);
not(t_344, d18);
not(t_345, o16);
and(c19, t_344, t_345);
not(t_346, o17);
not(t_347, e18);
and(d19, t_346, t_347);
not(t_348, e18);
not(t_349, r16);
and(e19, t_348, t_349);
not(t_350, p17);
not(t_351, f18);
and(f19, t_350, t_351);
not(t_352, f18);
not(t_353, u16);
and(g19, t_352, t_353);
not(t_354, q17);
not(t_355, g18);
and(h19, t_354, t_355);
not(t_356, g18);
not(t_357, x16);
and(i19, t_356, t_357);
not(t_358, r17);
not(t_359, h18);
and(j19, t_358, t_359);
not(t_360, h18);
not(t_361, a17);
and(k19, t_360, t_361);
not(t_362, j18);
not(t_363, k18);
and(l19, t_362, t_363);
not(t_364, i18);
not(t_365, v3);
and(m19, t_364, t_365);
not(t_366, l18);
not(t_367, m18);
and(n19, t_366, t_367);
not(t_368, n18);
not(t_369, o18);
and(o19, t_368, t_369);
not(t_370, p18);
not(t_371, q18);
and(p19, t_370, t_371);
not(t_372, r18);
not(t_373, s18);
and(q19, t_372, t_373);
not(t_374, t18);
not(t_375, u18);
and(r19, t_374, t_375);
not(t_376, v18);
not(t_377, w18);
and(s19, t_376, t_377);
not(t_378, x18);
not(t_379, y18);
and(t19, t_378, t_379);
not(t_380, z18);
not(t_381, a19);
and(u19, t_380, t_381);
not(t_382, b19);
not(t_383, c19);
and(v19, t_382, t_383);
not(t_384, d19);
not(t_385, e19);
and(w19, t_384, t_385);
not(t_386, f19);
not(t_387, g19);
and(x19, t_386, t_387);
not(t_388, h19);
not(t_389, i19);
and(y19, t_388, t_389);
not(t_390, j19);
not(t_391, k19);
and(z19, t_390, t_391);
not(t_392, d17);
not(t_393, m19);
and(a20, t_392, t_393);
not(t_394, i18);
not(t_395, m19);
and(b20, t_394, t_395);
not(t_396, m19);
not(t_397, v3);
and(c20, t_396, t_397);
not(t_398, l19);
not(t_399, l4);
and(d20, t_398, t_399);
not(t_400, n19);
not(t_401, b5);
and(e20, t_400, t_401);
not(t_402, o19);
not(t_403, r5);
and(f20, t_402, t_403);
not(t_404, p19);
not(t_405, h6);
and(g20, t_404, t_405);
not(t_406, q19);
not(t_407, x6);
and(h20, t_406, t_407);
not(t_408, r19);
not(t_409, n7);
and(i20, t_408, t_409);
not(t_410, s19);
not(t_411, d8);
and(j20, t_410, t_411);
not(t_412, t19);
not(t_413, t8);
and(k20, t_412, t_413);
not(t_414, u19);
not(t_415, j9);
and(l20, t_414, t_415);
not(t_416, v19);
not(t_417, z9);
and(m20, t_416, t_417);
not(t_418, w19);
not(t_419, p10);
and(n20, t_418, t_419);
not(t_420, x19);
not(t_421, f11);
and(o20, t_420, t_421);
not(t_422, y19);
not(t_423, v11);
and(p20, t_422, t_423);
not(t_424, z19);
not(t_425, l12);
and(q20, t_424, t_425);
not(t_426, f3);
not(t_427, a20);
and(r20, t_426, t_427);
not(t_428, b20);
not(t_429, c20);
and(s20, t_428, t_429);
not(t_430, l19);
not(t_431, d20);
and(t20, t_430, t_431);
not(t_432, u17);
not(t_433, d20);
and(u20, t_432, t_433);
not(t_434, n19);
not(t_435, e20);
and(v20, t_434, t_435);
not(t_436, d20);
not(t_437, l4);
and(w20, t_436, t_437);
not(t_438, v17);
not(t_439, e20);
and(x20, t_438, t_439);
not(t_440, o19);
not(t_441, f20);
and(y20, t_440, t_441);
not(t_442, e20);
not(t_443, b5);
and(z20, t_442, t_443);
not(t_444, w17);
not(t_445, f20);
and(a21, t_444, t_445);
not(t_446, p19);
not(t_447, g20);
and(b21, t_446, t_447);
not(t_448, f20);
not(t_449, r5);
and(c21, t_448, t_449);
not(t_450, x17);
not(t_451, g20);
and(d21, t_450, t_451);
not(t_452, q19);
not(t_453, h20);
and(e21, t_452, t_453);
not(t_454, g20);
not(t_455, h6);
and(f21, t_454, t_455);
not(t_456, y17);
not(t_457, h20);
and(g21, t_456, t_457);
not(t_458, r19);
not(t_459, i20);
and(h21, t_458, t_459);
not(t_460, h20);
not(t_461, x6);
and(i21, t_460, t_461);
not(t_462, z17);
not(t_463, i20);
and(j21, t_462, t_463);
not(t_464, s19);
not(t_465, j20);
and(k21, t_464, t_465);
not(t_466, i20);
not(t_467, n7);
and(l21, t_466, t_467);
not(t_468, a18);
not(t_469, j20);
and(m21, t_468, t_469);
not(t_470, t19);
not(t_471, k20);
and(n21, t_470, t_471);
not(t_472, j20);
not(t_473, d8);
and(o21, t_472, t_473);
not(t_474, b18);
not(t_475, k20);
and(p21, t_474, t_475);
not(t_476, u19);
not(t_477, l20);
and(q21, t_476, t_477);
not(t_478, k20);
not(t_479, t8);
and(r21, t_478, t_479);
not(t_480, c18);
not(t_481, l20);
and(s21, t_480, t_481);
not(t_482, v19);
not(t_483, m20);
and(t21, t_482, t_483);
not(t_484, l20);
not(t_485, j9);
and(u21, t_484, t_485);
not(t_486, d18);
not(t_487, m20);
and(v21, t_486, t_487);
not(t_488, w19);
not(t_489, n20);
and(w21, t_488, t_489);
not(t_490, m20);
not(t_491, z9);
and(x21, t_490, t_491);
not(t_492, e18);
not(t_493, n20);
and(y21, t_492, t_493);
not(t_494, x19);
not(t_495, o20);
and(z21, t_494, t_495);
not(t_496, n20);
not(t_497, p10);
and(a22, t_496, t_497);
not(t_498, f18);
not(t_499, o20);
and(b22, t_498, t_499);
not(t_500, y19);
not(t_501, p20);
and(c22, t_500, t_501);
not(t_502, o20);
not(t_503, f11);
and(d22, t_502, t_503);
not(t_504, g18);
not(t_505, p20);
and(e22, t_504, t_505);
not(t_506, z19);
not(t_507, q20);
and(f22, t_506, t_507);
not(t_508, p20);
not(t_509, v11);
and(g22, t_508, t_509);
not(t_510, h18);
not(t_511, q20);
and(h22, t_510, t_511);
not(t_512, q20);
not(t_513, l12);
and(i22, t_512, t_513);
not(t_514, f3);
not(t_515, r20);
and(j22, t_514, t_515);
not(t_516, r20);
not(t_517, a20);
and(k22, t_516, t_517);
not(t_518, s20);
not(t_519, u20);
and(l22, t_518, t_519);
not(t_520, t20);
not(t_521, w20);
and(m22, t_520, t_521);
not(t_522, v20);
not(t_523, z20);
and(n22, t_522, t_523);
not(t_524, y20);
not(t_525, c21);
and(o22, t_524, t_525);
not(t_526, b21);
not(t_527, f21);
and(p22, t_526, t_527);
not(t_528, e21);
not(t_529, i21);
and(q22, t_528, t_529);
not(t_530, h21);
not(t_531, l21);
and(r22, t_530, t_531);
not(t_532, k21);
not(t_533, o21);
and(s22, t_532, t_533);
not(t_534, n21);
not(t_535, r21);
and(t22, t_534, t_535);
not(t_536, q21);
not(t_537, u21);
and(u22, t_536, t_537);
not(t_538, t21);
not(t_539, x21);
and(v22, t_538, t_539);
not(t_540, w21);
not(t_541, a22);
and(w22, t_540, t_541);
not(t_542, z21);
not(t_543, d22);
and(x22, t_542, t_543);
not(t_544, c22);
not(t_545, g22);
and(y22, t_544, t_545);
not(t_546, j22);
not(t_547, k22);
and(z22, t_546, t_547);
not(t_548, s20);
not(t_549, l22);
and(a23, t_548, t_549);
not(t_550, l22);
not(t_551, u20);
and(b23, t_550, t_551);
not(t_552, m22);
not(t_553, x20);
and(c23, t_552, t_553);
not(t_554, n22);
not(t_555, a21);
and(d23, t_554, t_555);
not(t_556, o22);
not(t_557, d21);
and(e23, t_556, t_557);
not(t_558, p22);
not(t_559, g21);
and(f23, t_558, t_559);
not(t_560, q22);
not(t_561, j21);
and(g23, t_560, t_561);
not(t_562, r22);
not(t_563, m21);
and(h23, t_562, t_563);
not(t_564, s22);
not(t_565, p21);
and(i23, t_564, t_565);
not(t_566, t22);
not(t_567, s21);
and(j23, t_566, t_567);
not(t_568, u22);
not(t_569, v21);
and(k23, t_568, t_569);
not(t_570, v22);
not(t_571, y21);
and(l23, t_570, t_571);
not(t_572, w22);
not(t_573, b22);
and(m23, t_572, t_573);
not(t_574, x22);
not(t_575, e22);
and(n23, t_574, t_575);
not(t_576, y22);
not(t_577, h22);
and(o23, t_576, t_577);
not(t_578, a23);
not(t_579, b23);
and(p23, t_578, t_579);
not(t_580, m22);
not(t_581, c23);
and(q23, t_580, t_581);
not(t_582, z22);
not(t_583, u3);
and(r23, t_582, t_583);
not(t_584, n22);
not(t_585, d23);
and(s23, t_584, t_585);
not(t_586, c23);
not(t_587, x20);
and(t23, t_586, t_587);
not(t_588, o22);
not(t_589, e23);
and(u23, t_588, t_589);
not(t_590, d23);
not(t_591, a21);
and(v23, t_590, t_591);
not(t_592, p22);
not(t_593, f23);
and(w23, t_592, t_593);
not(t_594, e23);
not(t_595, d21);
and(x23, t_594, t_595);
not(t_596, q22);
not(t_597, g23);
and(y23, t_596, t_597);
not(t_598, f23);
not(t_599, g21);
and(z23, t_598, t_599);
not(t_600, r22);
not(t_601, h23);
and(a24, t_600, t_601);
not(t_602, g23);
not(t_603, j21);
and(b24, t_602, t_603);
not(t_604, s22);
not(t_605, i23);
and(c24, t_604, t_605);
not(t_606, h23);
not(t_607, m21);
and(d24, t_606, t_607);
not(t_608, t22);
not(t_609, j23);
and(e24, t_608, t_609);
not(t_610, i23);
not(t_611, p21);
and(f24, t_610, t_611);
not(t_612, u22);
not(t_613, k23);
and(g24, t_612, t_613);
not(t_614, j23);
not(t_615, s21);
and(h24, t_614, t_615);
not(t_616, v22);
not(t_617, l23);
and(i24, t_616, t_617);
not(t_618, k23);
not(t_619, v21);
and(j24, t_618, t_619);
not(t_620, w22);
not(t_621, m23);
and(k24, t_620, t_621);
not(t_622, l23);
not(t_623, y21);
and(l24, t_622, t_623);
not(t_624, x22);
not(t_625, n23);
and(m24, t_624, t_625);
not(t_626, m23);
not(t_627, b22);
and(n24, t_626, t_627);
not(t_628, y22);
not(t_629, o23);
and(o24, t_628, t_629);
not(t_630, n23);
not(t_631, e22);
and(p24, t_630, t_631);
not(t_632, o23);
not(t_633, h22);
and(q24, t_632, t_633);
not(t_634, r20);
not(t_635, r23);
and(r24, t_634, t_635);
not(t_636, z22);
not(t_637, r23);
and(s24, t_636, t_637);
not(t_638, q23);
not(t_639, t23);
and(t24, t_638, t_639);
not(t_640, r23);
not(t_641, u3);
and(u24, t_640, t_641);
not(t_642, s23);
not(t_643, v23);
and(v24, t_642, t_643);
not(t_644, p23);
not(t_645, k4);
and(w24, t_644, t_645);
not(t_646, u23);
not(t_647, x23);
and(x24, t_646, t_647);
not(t_648, w23);
not(t_649, z23);
and(y24, t_648, t_649);
not(t_650, y23);
not(t_651, b24);
and(z24, t_650, t_651);
not(t_652, a24);
not(t_653, d24);
and(a25, t_652, t_653);
not(t_654, c24);
not(t_655, f24);
and(b25, t_654, t_655);
not(t_656, e24);
not(t_657, h24);
and(c25, t_656, t_657);
not(t_658, g24);
not(t_659, j24);
and(d25, t_658, t_659);
not(t_660, i24);
not(t_661, l24);
and(e25, t_660, t_661);
not(t_662, k24);
not(t_663, n24);
and(f25, t_662, t_663);
not(t_664, m24);
not(t_665, p24);
and(g25, t_664, t_665);
not(t_666, o24);
not(t_667, q24);
and(h25, t_666, t_667);
not(t_668, e3);
not(t_669, r24);
and(i25, t_668, t_669);
not(t_670, s24);
not(t_671, u24);
and(j25, t_670, t_671);
not(t_672, l22);
not(t_673, w24);
and(k25, t_672, t_673);
not(t_674, p23);
not(t_675, w24);
and(l25, t_674, t_675);
not(t_676, w24);
not(t_677, k4);
and(m25, t_676, t_677);
not(t_678, t24);
not(t_679, a5);
and(n25, t_678, t_679);
not(t_680, v24);
not(t_681, q5);
and(o25, t_680, t_681);
not(t_682, x24);
not(t_683, g6);
and(p25, t_682, t_683);
not(t_684, y24);
not(t_685, w6);
and(q25, t_684, t_685);
not(t_686, z24);
not(t_687, m7);
and(r25, t_686, t_687);
not(t_688, a25);
not(t_689, c8);
and(s25, t_688, t_689);
not(t_690, b25);
not(t_691, s8);
and(t25, t_690, t_691);
not(t_692, c25);
not(t_693, i9);
and(u25, t_692, t_693);
not(t_694, d25);
not(t_695, y9);
and(v25, t_694, t_695);
not(t_696, e25);
not(t_697, o10);
and(w25, t_696, t_697);
not(t_698, f25);
not(t_699, e11);
and(x25, t_698, t_699);
not(t_700, g25);
not(t_701, u11);
and(y25, t_700, t_701);
not(t_702, h25);
not(t_703, k12);
and(z25, t_702, t_703);
not(t_704, e3);
not(t_705, i25);
and(a26, t_704, t_705);
not(t_706, i25);
not(t_707, r24);
and(b26, t_706, t_707);
not(t_708, j25);
not(t_709, k25);
and(c26, t_708, t_709);
not(t_710, l25);
not(t_711, m25);
and(d26, t_710, t_711);
not(t_712, t24);
not(t_713, n25);
and(e26, t_712, t_713);
not(t_714, v24);
not(t_715, o25);
and(f26, t_714, t_715);
not(t_716, c23);
not(t_717, n25);
and(g26, t_716, t_717);
not(t_718, x24);
not(t_719, p25);
and(h26, t_718, t_719);
not(t_720, n25);
not(t_721, a5);
and(i26, t_720, t_721);
not(t_722, d23);
not(t_723, o25);
and(j26, t_722, t_723);
not(t_724, y24);
not(t_725, q25);
and(k26, t_724, t_725);
not(t_726, o25);
not(t_727, q5);
and(l26, t_726, t_727);
not(t_728, e23);
not(t_729, p25);
and(m26, t_728, t_729);
not(t_730, z24);
not(t_731, r25);
and(n26, t_730, t_731);
not(t_732, p25);
not(t_733, g6);
and(o26, t_732, t_733);
not(t_734, f23);
not(t_735, q25);
and(p26, t_734, t_735);
not(t_736, a25);
not(t_737, s25);
and(q26, t_736, t_737);
not(t_738, q25);
not(t_739, w6);
and(r26, t_738, t_739);
not(t_740, g23);
not(t_741, r25);
and(s26, t_740, t_741);
not(t_742, b25);
not(t_743, t25);
and(t26, t_742, t_743);
not(t_744, r25);
not(t_745, m7);
and(u26, t_744, t_745);
not(t_746, h23);
not(t_747, s25);
and(v26, t_746, t_747);
not(t_748, c25);
not(t_749, u25);
and(w26, t_748, t_749);
not(t_750, s25);
not(t_751, c8);
and(x26, t_750, t_751);
not(t_752, i23);
not(t_753, t25);
and(y26, t_752, t_753);
not(t_754, d25);
not(t_755, v25);
and(z26, t_754, t_755);
not(t_756, t25);
not(t_757, s8);
and(a27, t_756, t_757);
not(t_758, j23);
not(t_759, u25);
and(b27, t_758, t_759);
not(t_760, e25);
not(t_761, w25);
and(c27, t_760, t_761);
not(t_762, u25);
not(t_763, i9);
and(d27, t_762, t_763);
not(t_764, k23);
not(t_765, v25);
and(e27, t_764, t_765);
not(t_766, f25);
not(t_767, x25);
and(f27, t_766, t_767);
not(t_768, v25);
not(t_769, y9);
and(g27, t_768, t_769);
not(t_770, l23);
not(t_771, w25);
and(h27, t_770, t_771);
not(t_772, g25);
not(t_773, y25);
and(i27, t_772, t_773);
not(t_774, w25);
not(t_775, o10);
and(j27, t_774, t_775);
not(t_776, m23);
not(t_777, x25);
and(k27, t_776, t_777);
not(t_778, h25);
not(t_779, z25);
and(l27, t_778, t_779);
not(t_780, x25);
not(t_781, e11);
and(m27, t_780, t_781);
not(t_782, n23);
not(t_783, y25);
and(n27, t_782, t_783);
not(t_784, y25);
not(t_785, u11);
and(o27, t_784, t_785);
not(t_786, o23);
not(t_787, z25);
and(p27, t_786, t_787);
not(t_788, z25);
not(t_789, k12);
and(q27, t_788, t_789);
not(t_790, a26);
not(t_791, b26);
and(r27, t_790, t_791);
not(t_792, j25);
not(t_793, c26);
and(s27, t_792, t_793);
not(t_794, c26);
not(t_795, k25);
and(t27, t_794, t_795);
not(t_796, d26);
not(t_797, g26);
and(u27, t_796, t_797);
not(t_798, e26);
not(t_799, i26);
and(v27, t_798, t_799);
not(t_800, f26);
not(t_801, l26);
and(w27, t_800, t_801);
not(t_802, h26);
not(t_803, o26);
and(x27, t_802, t_803);
not(t_804, k26);
not(t_805, r26);
and(y27, t_804, t_805);
not(t_806, n26);
not(t_807, u26);
and(z27, t_806, t_807);
not(t_808, q26);
not(t_809, x26);
and(a28, t_808, t_809);
not(t_810, t26);
not(t_811, a27);
and(b28, t_810, t_811);
not(t_812, w26);
not(t_813, d27);
and(c28, t_812, t_813);
not(t_814, z26);
not(t_815, g27);
and(d28, t_814, t_815);
not(t_816, c27);
not(t_817, j27);
and(e28, t_816, t_817);
not(t_818, f27);
not(t_819, m27);
and(f28, t_818, t_819);
not(t_820, i27);
not(t_821, o27);
and(g28, t_820, t_821);
not(t_822, s27);
not(t_823, t27);
and(h28, t_822, t_823);
not(t_824, d26);
not(t_825, u27);
and(i28, t_824, t_825);
not(t_826, r27);
not(t_827, t3);
and(j28, t_826, t_827);
not(t_828, u27);
not(t_829, g26);
and(k28, t_828, t_829);
not(t_830, v27);
not(t_831, j26);
and(l28, t_830, t_831);
not(t_832, w27);
not(t_833, m26);
and(m28, t_832, t_833);
not(t_834, x27);
not(t_835, p26);
and(n28, t_834, t_835);
not(t_836, y27);
not(t_837, s26);
and(o28, t_836, t_837);
not(t_838, z27);
not(t_839, v26);
and(p28, t_838, t_839);
not(t_840, a28);
not(t_841, y26);
and(q28, t_840, t_841);
not(t_842, b28);
not(t_843, b27);
and(r28, t_842, t_843);
not(t_844, c28);
not(t_845, e27);
and(s28, t_844, t_845);
not(t_846, d28);
not(t_847, h27);
and(t28, t_846, t_847);
not(t_848, e28);
not(t_849, k27);
and(u28, t_848, t_849);
not(t_850, f28);
not(t_851, n27);
and(v28, t_850, t_851);
not(t_852, g28);
not(t_853, p27);
and(w28, t_852, t_853);
not(t_854, i25);
not(t_855, j28);
and(x28, t_854, t_855);
not(t_856, r27);
not(t_857, j28);
and(y28, t_856, t_857);
not(t_858, i28);
not(t_859, k28);
and(z28, t_858, t_859);
not(t_860, v27);
not(t_861, l28);
and(a29, t_860, t_861);
not(t_862, j28);
not(t_863, t3);
and(b29, t_862, t_863);
not(t_864, w27);
not(t_865, m28);
and(c29, t_864, t_865);
not(t_866, h28);
not(t_867, j4);
and(d29, t_866, t_867);
not(t_868, x27);
not(t_869, n28);
and(e29, t_868, t_869);
not(t_870, l28);
not(t_871, j26);
and(f29, t_870, t_871);
not(t_872, y27);
not(t_873, o28);
and(g29, t_872, t_873);
not(t_874, m28);
not(t_875, m26);
and(h29, t_874, t_875);
not(t_876, z27);
not(t_877, p28);
and(i29, t_876, t_877);
not(t_878, n28);
not(t_879, p26);
and(j29, t_878, t_879);
not(t_880, a28);
not(t_881, q28);
and(k29, t_880, t_881);
not(t_882, o28);
not(t_883, s26);
and(l29, t_882, t_883);
not(t_884, b28);
not(t_885, r28);
and(m29, t_884, t_885);
not(t_886, p28);
not(t_887, v26);
and(n29, t_886, t_887);
not(t_888, c28);
not(t_889, s28);
and(o29, t_888, t_889);
not(t_890, q28);
not(t_891, y26);
and(p29, t_890, t_891);
not(t_892, d28);
not(t_893, t28);
and(q29, t_892, t_893);
not(t_894, r28);
not(t_895, b27);
and(r29, t_894, t_895);
not(t_896, e28);
not(t_897, u28);
and(s29, t_896, t_897);
not(t_898, s28);
not(t_899, e27);
and(t29, t_898, t_899);
not(t_900, f28);
not(t_901, v28);
and(u29, t_900, t_901);
not(t_902, t28);
not(t_903, h27);
and(v29, t_902, t_903);
not(t_904, g28);
not(t_905, w28);
and(w29, t_904, t_905);
not(t_906, u28);
not(t_907, k27);
and(x29, t_906, t_907);
not(t_908, v28);
not(t_909, n27);
and(y29, t_908, t_909);
not(t_910, w28);
not(t_911, p27);
and(z29, t_910, t_911);
not(t_912, d3);
not(t_913, x28);
and(a30, t_912, t_913);
not(t_914, y28);
not(t_915, b29);
and(b30, t_914, t_915);
not(t_916, c26);
not(t_917, d29);
and(c30, t_916, t_917);
not(t_918, h28);
not(t_919, d29);
and(d30, t_918, t_919);
not(t_920, a29);
not(t_921, f29);
and(e30, t_920, t_921);
not(t_922, c29);
not(t_923, h29);
and(f30, t_922, t_923);
not(t_924, d29);
not(t_925, j4);
and(g30, t_924, t_925);
not(t_926, e29);
not(t_927, j29);
and(h30, t_926, t_927);
not(t_928, z28);
not(t_929, z4);
and(i30, t_928, t_929);
not(t_930, g29);
not(t_931, l29);
and(j30, t_930, t_931);
not(t_932, i29);
not(t_933, n29);
and(k30, t_932, t_933);
not(t_934, k29);
not(t_935, p29);
and(l30, t_934, t_935);
not(t_936, m29);
not(t_937, r29);
and(m30, t_936, t_937);
not(t_938, o29);
not(t_939, t29);
and(n30, t_938, t_939);
not(t_940, q29);
not(t_941, v29);
and(o30, t_940, t_941);
not(t_942, s29);
not(t_943, x29);
and(p30, t_942, t_943);
not(t_944, u29);
not(t_945, y29);
and(q30, t_944, t_945);
not(t_946, w29);
not(t_947, z29);
and(r30, t_946, t_947);
not(t_948, d3);
not(t_949, a30);
and(s30, t_948, t_949);
not(t_950, a30);
not(t_951, x28);
and(t30, t_950, t_951);
not(t_952, b30);
not(t_953, c30);
and(u30, t_952, t_953);
not(t_954, d30);
not(t_955, g30);
and(v30, t_954, t_955);
not(t_956, u27);
not(t_957, i30);
and(w30, t_956, t_957);
not(t_958, z28);
not(t_959, i30);
and(x30, t_958, t_959);
not(t_960, i30);
not(t_961, z4);
and(y30, t_960, t_961);
not(t_962, e30);
not(t_963, p5);
and(z30, t_962, t_963);
not(t_964, f30);
not(t_965, f6);
and(a31, t_964, t_965);
not(t_966, h30);
not(t_967, v6);
and(b31, t_966, t_967);
not(t_968, j30);
not(t_969, l7);
and(c31, t_968, t_969);
not(t_970, k30);
not(t_971, b8);
and(d31, t_970, t_971);
not(t_972, l30);
not(t_973, r8);
and(e31, t_972, t_973);
not(t_974, m30);
not(t_975, h9);
and(f31, t_974, t_975);
not(t_976, n30);
not(t_977, x9);
and(g31, t_976, t_977);
not(t_978, o30);
not(t_979, n10);
and(h31, t_978, t_979);
not(t_980, p30);
not(t_981, d11);
and(i31, t_980, t_981);
not(t_982, q30);
not(t_983, t11);
and(j31, t_982, t_983);
not(t_984, r30);
not(t_985, j12);
and(k31, t_984, t_985);
not(t_986, s30);
not(t_987, t30);
and(l31, t_986, t_987);
not(t_988, b30);
not(t_989, u30);
and(m31, t_988, t_989);
not(t_990, u30);
not(t_991, c30);
and(n31, t_990, t_991);
not(t_992, v30);
not(t_993, w30);
and(o31, t_992, t_993);
not(t_994, x30);
not(t_995, y30);
and(p31, t_994, t_995);
not(t_996, e30);
not(t_997, z30);
and(q31, t_996, t_997);
not(t_998, f30);
not(t_999, a31);
and(r31, t_998, t_999);
not(t_1000, h30);
not(t_1001, b31);
and(s31, t_1000, t_1001);
not(t_1002, l28);
not(t_1003, z30);
and(t31, t_1002, t_1003);
not(t_1004, j30);
not(t_1005, c31);
and(u31, t_1004, t_1005);
not(t_1006, z30);
not(t_1007, p5);
and(v31, t_1006, t_1007);
not(t_1008, m28);
not(t_1009, a31);
and(w31, t_1008, t_1009);
not(t_1010, k30);
not(t_1011, d31);
and(x31, t_1010, t_1011);
not(t_1012, a31);
not(t_1013, f6);
and(y31, t_1012, t_1013);
not(t_1014, n28);
not(t_1015, b31);
and(z31, t_1014, t_1015);
not(t_1016, l30);
not(t_1017, e31);
and(a32, t_1016, t_1017);
not(t_1018, b31);
not(t_1019, v6);
and(b32, t_1018, t_1019);
not(t_1020, o28);
not(t_1021, c31);
and(c32, t_1020, t_1021);
not(t_1022, m30);
not(t_1023, f31);
and(d32, t_1022, t_1023);
not(t_1024, c31);
not(t_1025, l7);
and(e32, t_1024, t_1025);
not(t_1026, p28);
not(t_1027, d31);
and(f32, t_1026, t_1027);
not(t_1028, n30);
not(t_1029, g31);
and(g32, t_1028, t_1029);
not(t_1030, d31);
not(t_1031, b8);
and(h32, t_1030, t_1031);
not(t_1032, q28);
not(t_1033, e31);
and(i32, t_1032, t_1033);
not(t_1034, o30);
not(t_1035, h31);
and(j32, t_1034, t_1035);
not(t_1036, e31);
not(t_1037, r8);
and(k32, t_1036, t_1037);
not(t_1038, r28);
not(t_1039, f31);
and(l32, t_1038, t_1039);
not(t_1040, p30);
not(t_1041, i31);
and(m32, t_1040, t_1041);
not(t_1042, f31);
not(t_1043, h9);
and(n32, t_1042, t_1043);
not(t_1044, s28);
not(t_1045, g31);
and(o32, t_1044, t_1045);
not(t_1046, q30);
not(t_1047, j31);
and(p32, t_1046, t_1047);
not(t_1048, g31);
not(t_1049, x9);
and(q32, t_1048, t_1049);
not(t_1050, t28);
not(t_1051, h31);
and(r32, t_1050, t_1051);
not(t_1052, r30);
not(t_1053, k31);
and(s32, t_1052, t_1053);
not(t_1054, h31);
not(t_1055, n10);
and(t32, t_1054, t_1055);
not(t_1056, u28);
not(t_1057, i31);
and(u32, t_1056, t_1057);
not(t_1058, i31);
not(t_1059, d11);
and(v32, t_1058, t_1059);
not(t_1060, v28);
not(t_1061, j31);
and(w32, t_1060, t_1061);
not(t_1062, j31);
not(t_1063, t11);
and(x32, t_1062, t_1063);
not(t_1064, w28);
not(t_1065, k31);
and(y32, t_1064, t_1065);
not(t_1066, k31);
not(t_1067, j12);
and(z32, t_1066, t_1067);
not(t_1068, m31);
not(t_1069, n31);
and(a33, t_1068, t_1069);
not(t_1070, v30);
not(t_1071, o31);
and(b33, t_1070, t_1071);
not(t_1072, o31);
not(t_1073, w30);
and(c33, t_1072, t_1073);
not(t_1074, p31);
not(t_1075, t31);
and(d33, t_1074, t_1075);
not(t_1076, q31);
not(t_1077, v31);
and(e33, t_1076, t_1077);
not(t_1078, l31);
not(t_1079, s3);
and(f33, t_1078, t_1079);
not(t_1080, r31);
not(t_1081, y31);
and(g33, t_1080, t_1081);
not(t_1082, s31);
not(t_1083, b32);
and(h33, t_1082, t_1083);
not(t_1084, u31);
not(t_1085, e32);
and(i33, t_1084, t_1085);
not(t_1086, x31);
not(t_1087, h32);
and(j33, t_1086, t_1087);
not(t_1088, a32);
not(t_1089, k32);
and(k33, t_1088, t_1089);
not(t_1090, d32);
not(t_1091, n32);
and(l33, t_1090, t_1091);
not(t_1092, g32);
not(t_1093, q32);
and(m33, t_1092, t_1093);
not(t_1094, j32);
not(t_1095, t32);
and(n33, t_1094, t_1095);
not(t_1096, m32);
not(t_1097, v32);
and(o33, t_1096, t_1097);
not(t_1098, p32);
not(t_1099, x32);
and(p33, t_1098, t_1099);
not(t_1100, a30);
not(t_1101, f33);
and(q33, t_1100, t_1101);
not(t_1102, l31);
not(t_1103, f33);
and(r33, t_1102, t_1103);
not(t_1104, b33);
not(t_1105, c33);
and(s33, t_1104, t_1105);
not(t_1106, p31);
not(t_1107, d33);
and(t33, t_1106, t_1107);
not(t_1108, f33);
not(t_1109, s3);
and(u33, t_1108, t_1109);
not(t_1110, a33);
not(t_1111, i4);
and(v33, t_1110, t_1111);
not(t_1112, d33);
not(t_1113, t31);
and(w33, t_1112, t_1113);
not(t_1114, e33);
not(t_1115, w31);
and(x33, t_1114, t_1115);
not(t_1116, g33);
not(t_1117, z31);
and(y33, t_1116, t_1117);
not(t_1118, h33);
not(t_1119, c32);
and(z33, t_1118, t_1119);
not(t_1120, i33);
not(t_1121, f32);
and(a34, t_1120, t_1121);
not(t_1122, j33);
not(t_1123, i32);
and(b34, t_1122, t_1123);
not(t_1124, k33);
not(t_1125, l32);
and(c34, t_1124, t_1125);
not(t_1126, l33);
not(t_1127, o32);
and(d34, t_1126, t_1127);
not(t_1128, m33);
not(t_1129, r32);
and(e34, t_1128, t_1129);
not(t_1130, n33);
not(t_1131, u32);
and(f34, t_1130, t_1131);
not(t_1132, o33);
not(t_1133, w32);
and(g34, t_1132, t_1133);
not(t_1134, p33);
not(t_1135, y32);
and(h34, t_1134, t_1135);
not(t_1136, c3);
not(t_1137, q33);
and(i34, t_1136, t_1137);
not(t_1138, r33);
not(t_1139, u33);
and(j34, t_1138, t_1139);
not(t_1140, u30);
not(t_1141, v33);
and(k34, t_1140, t_1141);
not(t_1142, a33);
not(t_1143, v33);
and(l34, t_1142, t_1143);
not(t_1144, t33);
not(t_1145, w33);
and(m34, t_1144, t_1145);
not(t_1146, e33);
not(t_1147, x33);
and(n34, t_1146, t_1147);
not(t_1148, g33);
not(t_1149, y33);
and(o34, t_1148, t_1149);
not(t_1150, v33);
not(t_1151, i4);
and(p34, t_1150, t_1151);
not(t_1152, h33);
not(t_1153, z33);
and(q34, t_1152, t_1153);
not(t_1154, s33);
not(t_1155, y4);
and(r34, t_1154, t_1155);
not(t_1156, i33);
not(t_1157, a34);
and(s34, t_1156, t_1157);
not(t_1158, x33);
not(t_1159, w31);
and(t34, t_1158, t_1159);
not(t_1160, j33);
not(t_1161, b34);
and(u34, t_1160, t_1161);
not(t_1162, y33);
not(t_1163, z31);
and(v34, t_1162, t_1163);
not(t_1164, k33);
not(t_1165, c34);
and(w34, t_1164, t_1165);
not(t_1166, z33);
not(t_1167, c32);
and(x34, t_1166, t_1167);
not(t_1168, l33);
not(t_1169, d34);
and(y34, t_1168, t_1169);
not(t_1170, a34);
not(t_1171, f32);
and(z34, t_1170, t_1171);
not(t_1172, m33);
not(t_1173, e34);
and(a35, t_1172, t_1173);
not(t_1174, b34);
not(t_1175, i32);
and(b35, t_1174, t_1175);
not(t_1176, n33);
not(t_1177, f34);
and(c35, t_1176, t_1177);
not(t_1178, c34);
not(t_1179, l32);
and(d35, t_1178, t_1179);
not(t_1180, o33);
not(t_1181, g34);
and(e35, t_1180, t_1181);
not(t_1182, d34);
not(t_1183, o32);
and(f35, t_1182, t_1183);
not(t_1184, p33);
not(t_1185, h34);
and(g35, t_1184, t_1185);
not(t_1186, e34);
not(t_1187, r32);
and(h35, t_1186, t_1187);
not(t_1188, f34);
not(t_1189, u32);
and(i35, t_1188, t_1189);
not(t_1190, g34);
not(t_1191, w32);
and(j35, t_1190, t_1191);
not(t_1192, h34);
not(t_1193, y32);
and(k35, t_1192, t_1193);
not(t_1194, c3);
not(t_1195, i34);
and(l35, t_1194, t_1195);
not(t_1196, i34);
not(t_1197, q33);
and(m35, t_1196, t_1197);
not(t_1198, j34);
not(t_1199, k34);
and(n35, t_1198, t_1199);
not(t_1200, l34);
not(t_1201, p34);
and(o35, t_1200, t_1201);
not(t_1202, o31);
not(t_1203, r34);
and(p35, t_1202, t_1203);
not(t_1204, s33);
not(t_1205, r34);
and(q35, t_1204, t_1205);
not(t_1206, n34);
not(t_1207, t34);
and(r35, t_1206, t_1207);
not(t_1208, o34);
not(t_1209, v34);
and(s35, t_1208, t_1209);
not(t_1210, q34);
not(t_1211, x34);
and(t35, t_1210, t_1211);
not(t_1212, r34);
not(t_1213, y4);
and(u35, t_1212, t_1213);
not(t_1214, s34);
not(t_1215, z34);
and(v35, t_1214, t_1215);
not(t_1216, m34);
not(t_1217, o5);
and(w35, t_1216, t_1217);
not(t_1218, u34);
not(t_1219, b35);
and(x35, t_1218, t_1219);
not(t_1220, w34);
not(t_1221, d35);
and(y35, t_1220, t_1221);
not(t_1222, y34);
not(t_1223, f35);
and(z35, t_1222, t_1223);
not(t_1224, a35);
not(t_1225, h35);
and(a36, t_1224, t_1225);
not(t_1226, c35);
not(t_1227, i35);
and(b36, t_1226, t_1227);
not(t_1228, e35);
not(t_1229, j35);
and(c36, t_1228, t_1229);
not(t_1230, g35);
not(t_1231, k35);
and(d36, t_1230, t_1231);
not(t_1232, l35);
not(t_1233, m35);
and(e36, t_1232, t_1233);
not(t_1234, j34);
not(t_1235, n35);
and(f36, t_1234, t_1235);
not(t_1236, n35);
not(t_1237, k34);
and(g36, t_1236, t_1237);
not(t_1238, o35);
not(t_1239, p35);
and(h36, t_1238, t_1239);
not(t_1240, q35);
not(t_1241, u35);
and(i36, t_1240, t_1241);
not(t_1242, d33);
not(t_1243, w35);
and(j36, t_1242, t_1243);
not(t_1244, m34);
not(t_1245, w35);
and(k36, t_1244, t_1245);
not(t_1246, w35);
not(t_1247, o5);
and(l36, t_1246, t_1247);
not(t_1248, r35);
not(t_1249, e6);
and(m36, t_1248, t_1249);
not(t_1250, s35);
not(t_1251, u6);
and(n36, t_1250, t_1251);
not(t_1252, t35);
not(t_1253, k7);
and(o36, t_1252, t_1253);
not(t_1254, v35);
not(t_1255, a8);
and(p36, t_1254, t_1255);
not(t_1256, x35);
not(t_1257, q8);
and(q36, t_1256, t_1257);
not(t_1258, y35);
not(t_1259, g9);
and(r36, t_1258, t_1259);
not(t_1260, z35);
not(t_1261, w9);
and(s36, t_1260, t_1261);
not(t_1262, a36);
not(t_1263, m10);
and(t36, t_1262, t_1263);
not(t_1264, b36);
not(t_1265, c11);
and(u36, t_1264, t_1265);
not(t_1266, c36);
not(t_1267, s11);
and(v36, t_1266, t_1267);
not(t_1268, d36);
not(t_1269, i12);
and(w36, t_1268, t_1269);
not(t_1270, f36);
not(t_1271, g36);
and(x36, t_1270, t_1271);
not(t_1272, o35);
not(t_1273, h36);
and(y36, t_1272, t_1273);
not(t_1274, h36);
not(t_1275, p35);
and(z36, t_1274, t_1275);
not(t_1276, i36);
not(t_1277, j36);
and(a37, t_1276, t_1277);
not(t_1278, k36);
not(t_1279, l36);
and(b37, t_1278, t_1279);
not(t_1280, r35);
not(t_1281, m36);
and(c37, t_1280, t_1281);
not(t_1282, e36);
not(t_1283, r3);
and(d37, t_1282, t_1283);
not(t_1284, s35);
not(t_1285, n36);
and(e37, t_1284, t_1285);
not(t_1286, t35);
not(t_1287, o36);
and(f37, t_1286, t_1287);
not(t_1288, v35);
not(t_1289, p36);
and(g37, t_1288, t_1289);
not(t_1290, x33);
not(t_1291, m36);
and(h37, t_1290, t_1291);
not(t_1292, x35);
not(t_1293, q36);
and(i37, t_1292, t_1293);
not(t_1294, m36);
not(t_1295, e6);
and(j37, t_1294, t_1295);
not(t_1296, y33);
not(t_1297, n36);
and(k37, t_1296, t_1297);
not(t_1298, y35);
not(t_1299, r36);
and(l37, t_1298, t_1299);
not(t_1300, n36);
not(t_1301, u6);
and(m37, t_1300, t_1301);
not(t_1302, z33);
not(t_1303, o36);
and(n37, t_1302, t_1303);
not(t_1304, z35);
not(t_1305, s36);
and(o37, t_1304, t_1305);
not(t_1306, o36);
not(t_1307, k7);
and(p37, t_1306, t_1307);
not(t_1308, a34);
not(t_1309, p36);
and(q37, t_1308, t_1309);
not(t_1310, a36);
not(t_1311, t36);
and(r37, t_1310, t_1311);
not(t_1312, p36);
not(t_1313, a8);
and(s37, t_1312, t_1313);
not(t_1314, b34);
not(t_1315, q36);
and(t37, t_1314, t_1315);
not(t_1316, b36);
not(t_1317, u36);
and(u37, t_1316, t_1317);
not(t_1318, q36);
not(t_1319, q8);
and(v37, t_1318, t_1319);
not(t_1320, c34);
not(t_1321, r36);
and(w37, t_1320, t_1321);
not(t_1322, c36);
not(t_1323, v36);
and(x37, t_1322, t_1323);
not(t_1324, r36);
not(t_1325, g9);
and(y37, t_1324, t_1325);
not(t_1326, d34);
not(t_1327, s36);
and(z37, t_1326, t_1327);
not(t_1328, d36);
not(t_1329, w36);
and(a38, t_1328, t_1329);
not(t_1330, s36);
not(t_1331, w9);
and(b38, t_1330, t_1331);
not(t_1332, e34);
not(t_1333, t36);
and(c38, t_1332, t_1333);
not(t_1334, t36);
not(t_1335, m10);
and(d38, t_1334, t_1335);
not(t_1336, f34);
not(t_1337, u36);
and(e38, t_1336, t_1337);
not(t_1338, u36);
not(t_1339, c11);
and(f38, t_1338, t_1339);
not(t_1340, g34);
not(t_1341, v36);
and(g38, t_1340, t_1341);
not(t_1342, v36);
not(t_1343, s11);
and(h38, t_1342, t_1343);
not(t_1344, h34);
not(t_1345, w36);
and(i38, t_1344, t_1345);
not(t_1346, w36);
not(t_1347, i12);
and(j38, t_1346, t_1347);
not(t_1348, i34);
not(t_1349, d37);
and(k38, t_1348, t_1349);
not(t_1350, e36);
not(t_1351, d37);
and(l38, t_1350, t_1351);
not(t_1352, y36);
not(t_1353, z36);
and(m38, t_1352, t_1353);
not(t_1354, i36);
not(t_1355, a37);
and(n38, t_1354, t_1355);
not(t_1356, a37);
not(t_1357, j36);
and(o38, t_1356, t_1357);
not(t_1358, b37);
not(t_1359, h37);
and(p38, t_1358, t_1359);
not(t_1360, c37);
not(t_1361, j37);
and(q38, t_1360, t_1361);
not(t_1362, d37);
not(t_1363, r3);
and(r38, t_1362, t_1363);
not(t_1364, e37);
not(t_1365, m37);
and(s38, t_1364, t_1365);
not(t_1366, x36);
not(t_1367, h4);
and(t38, t_1366, t_1367);
not(t_1368, f37);
not(t_1369, p37);
and(u38, t_1368, t_1369);
not(t_1370, g37);
not(t_1371, s37);
and(v38, t_1370, t_1371);
not(t_1372, i37);
not(t_1373, v37);
and(w38, t_1372, t_1373);
not(t_1374, l37);
not(t_1375, y37);
and(x38, t_1374, t_1375);
not(t_1376, o37);
not(t_1377, b38);
and(y38, t_1376, t_1377);
not(t_1378, r37);
not(t_1379, d38);
and(z38, t_1378, t_1379);
not(t_1380, u37);
not(t_1381, f38);
and(a39, t_1380, t_1381);
not(t_1382, x37);
not(t_1383, h38);
and(b39, t_1382, t_1383);
not(t_1384, b3);
not(t_1385, k38);
and(c39, t_1384, t_1385);
not(t_1386, l38);
not(t_1387, r38);
and(d39, t_1386, t_1387);
not(t_1388, n35);
not(t_1389, t38);
and(e39, t_1388, t_1389);
not(t_1390, x36);
not(t_1391, t38);
and(f39, t_1390, t_1391);
not(t_1392, n38);
not(t_1393, o38);
and(g39, t_1392, t_1393);
not(t_1394, b37);
not(t_1395, p38);
and(h39, t_1394, t_1395);
not(t_1396, t38);
not(t_1397, h4);
and(i39, t_1396, t_1397);
not(t_1398, m38);
not(t_1399, x4);
and(j39, t_1398, t_1399);
not(t_1400, p38);
not(t_1401, h37);
and(k39, t_1400, t_1401);
not(t_1402, q38);
not(t_1403, k37);
and(l39, t_1402, t_1403);
not(t_1404, s38);
not(t_1405, n37);
and(m39, t_1404, t_1405);
not(t_1406, u38);
not(t_1407, q37);
and(n39, t_1406, t_1407);
not(t_1408, v38);
not(t_1409, t37);
and(o39, t_1408, t_1409);
not(t_1410, w38);
not(t_1411, w37);
and(p39, t_1410, t_1411);
not(t_1412, x38);
not(t_1413, z37);
and(q39, t_1412, t_1413);
not(t_1414, y38);
not(t_1415, c38);
and(r39, t_1414, t_1415);
not(t_1416, z38);
not(t_1417, e38);
and(s39, t_1416, t_1417);
not(t_1418, a39);
not(t_1419, g38);
and(t39, t_1418, t_1419);
not(t_1420, b39);
not(t_1421, i38);
and(u39, t_1420, t_1421);
not(t_1422, b3);
not(t_1423, c39);
and(v39, t_1422, t_1423);
not(t_1424, c39);
not(t_1425, k38);
and(w39, t_1424, t_1425);
not(t_1426, d39);
not(t_1427, e39);
and(x39, t_1426, t_1427);
not(t_1428, f39);
not(t_1429, i39);
and(y39, t_1428, t_1429);
not(t_1430, h36);
not(t_1431, j39);
and(z39, t_1430, t_1431);
not(t_1432, m38);
not(t_1433, j39);
and(a40, t_1432, t_1433);
not(t_1434, h39);
not(t_1435, k39);
and(b40, t_1434, t_1435);
not(t_1436, q38);
not(t_1437, l39);
and(c40, t_1436, t_1437);
not(t_1438, s38);
not(t_1439, m39);
and(d40, t_1438, t_1439);
not(t_1440, u38);
not(t_1441, n39);
and(e40, t_1440, t_1441);
not(t_1442, j39);
not(t_1443, x4);
and(f40, t_1442, t_1443);
not(t_1444, v38);
not(t_1445, o39);
and(g40, t_1444, t_1445);
not(t_1446, g39);
not(t_1447, n5);
and(h40, t_1446, t_1447);
not(t_1448, w38);
not(t_1449, p39);
and(i40, t_1448, t_1449);
not(t_1450, l39);
not(t_1451, k37);
and(j40, t_1450, t_1451);
not(t_1452, x38);
not(t_1453, q39);
and(k40, t_1452, t_1453);
not(t_1454, m39);
not(t_1455, n37);
and(l40, t_1454, t_1455);
not(t_1456, y38);
not(t_1457, r39);
and(m40, t_1456, t_1457);
not(t_1458, n39);
not(t_1459, q37);
and(n40, t_1458, t_1459);
not(t_1460, z38);
not(t_1461, s39);
and(o40, t_1460, t_1461);
not(t_1462, o39);
not(t_1463, t37);
and(p40, t_1462, t_1463);
not(t_1464, a39);
not(t_1465, t39);
and(q40, t_1464, t_1465);
not(t_1466, p39);
not(t_1467, w37);
and(r40, t_1466, t_1467);
not(t_1468, b39);
not(t_1469, u39);
and(s40, t_1468, t_1469);
not(t_1470, q39);
not(t_1471, z37);
and(t40, t_1470, t_1471);
not(t_1472, r39);
not(t_1473, c38);
and(u40, t_1472, t_1473);
not(t_1474, s39);
not(t_1475, e38);
and(v40, t_1474, t_1475);
not(t_1476, t39);
not(t_1477, g38);
and(w40, t_1476, t_1477);
not(t_1478, u39);
not(t_1479, i38);
and(x40, t_1478, t_1479);
not(t_1480, v39);
not(t_1481, w39);
and(y40, t_1480, t_1481);
not(t_1482, d39);
not(t_1483, x39);
and(z40, t_1482, t_1483);
not(t_1484, x39);
not(t_1485, e39);
and(a41, t_1484, t_1485);
not(t_1486, y39);
not(t_1487, z39);
and(b41, t_1486, t_1487);
not(t_1488, a40);
not(t_1489, f40);
and(c41, t_1488, t_1489);
not(t_1490, a37);
not(t_1491, h40);
and(d41, t_1490, t_1491);
not(t_1492, g39);
not(t_1493, h40);
and(e41, t_1492, t_1493);
not(t_1494, c40);
not(t_1495, j40);
and(f41, t_1494, t_1495);
not(t_1496, d40);
not(t_1497, l40);
and(g41, t_1496, t_1497);
not(t_1498, e40);
not(t_1499, n40);
and(h41, t_1498, t_1499);
not(t_1500, g40);
not(t_1501, p40);
and(i41, t_1500, t_1501);
not(t_1502, h40);
not(t_1503, n5);
and(j41, t_1502, t_1503);
not(t_1504, i40);
not(t_1505, r40);
and(k41, t_1504, t_1505);
not(t_1506, b40);
not(t_1507, d6);
and(l41, t_1506, t_1507);
not(t_1508, k40);
not(t_1509, t40);
and(m41, t_1508, t_1509);
not(t_1510, m40);
not(t_1511, u40);
and(n41, t_1510, t_1511);
not(t_1512, o40);
not(t_1513, v40);
and(o41, t_1512, t_1513);
not(t_1514, q40);
not(t_1515, w40);
and(p41, t_1514, t_1515);
not(t_1516, s40);
not(t_1517, x40);
and(q41, t_1516, t_1517);
not(t_1518, z40);
not(t_1519, a41);
and(r41, t_1518, t_1519);
not(t_1520, y39);
not(t_1521, b41);
and(s41, t_1520, t_1521);
not(t_1522, b41);
not(t_1523, z39);
and(t41, t_1522, t_1523);
not(t_1524, c41);
not(t_1525, d41);
and(u41, t_1524, t_1525);
not(t_1526, e41);
not(t_1527, j41);
and(v41, t_1526, t_1527);
not(t_1528, p38);
not(t_1529, l41);
and(w41, t_1528, t_1529);
not(t_1530, b40);
not(t_1531, l41);
and(x41, t_1530, t_1531);
not(t_1532, y40);
not(t_1533, q3);
and(y41, t_1532, t_1533);
not(t_1534, l41);
not(t_1535, d6);
and(z41, t_1534, t_1535);
not(t_1536, f41);
not(t_1537, t6);
and(a42, t_1536, t_1537);
not(t_1538, g41);
not(t_1539, j7);
and(b42, t_1538, t_1539);
not(t_1540, h41);
not(t_1541, z7);
and(c42, t_1540, t_1541);
not(t_1542, i41);
not(t_1543, p8);
and(d42, t_1542, t_1543);
not(t_1544, k41);
not(t_1545, f9);
and(e42, t_1544, t_1545);
not(t_1546, m41);
not(t_1547, v9);
and(f42, t_1546, t_1547);
not(t_1548, n41);
not(t_1549, l10);
and(g42, t_1548, t_1549);
not(t_1550, o41);
not(t_1551, b11);
and(h42, t_1550, t_1551);
not(t_1552, p41);
not(t_1553, r11);
and(i42, t_1552, t_1553);
not(t_1554, q41);
not(t_1555, h12);
and(j42, t_1554, t_1555);
not(t_1556, c39);
not(t_1557, y41);
and(k42, t_1556, t_1557);
not(t_1558, y40);
not(t_1559, y41);
and(l42, t_1558, t_1559);
not(t_1560, s41);
not(t_1561, t41);
and(m42, t_1560, t_1561);
not(t_1562, c41);
not(t_1563, u41);
and(n42, t_1562, t_1563);
not(t_1564, u41);
not(t_1565, d41);
and(o42, t_1564, t_1565);
not(t_1566, v41);
not(t_1567, w41);
and(p42, t_1566, t_1567);
not(t_1568, x41);
not(t_1569, z41);
and(q42, t_1568, t_1569);
not(t_1570, f41);
not(t_1571, a42);
and(r42, t_1570, t_1571);
not(t_1572, y41);
not(t_1573, q3);
and(s42, t_1572, t_1573);
not(t_1574, g41);
not(t_1575, b42);
and(t42, t_1574, t_1575);
not(t_1576, r41);
not(t_1577, g4);
and(u42, t_1576, t_1577);
not(t_1578, h41);
not(t_1579, c42);
and(v42, t_1578, t_1579);
not(t_1580, i41);
not(t_1581, d42);
and(w42, t_1580, t_1581);
not(t_1582, k41);
not(t_1583, e42);
and(x42, t_1582, t_1583);
not(t_1584, l39);
not(t_1585, a42);
and(y42, t_1584, t_1585);
not(t_1586, m41);
not(t_1587, f42);
and(z42, t_1586, t_1587);
not(t_1588, a42);
not(t_1589, t6);
and(a43, t_1588, t_1589);
not(t_1590, m39);
not(t_1591, b42);
and(b43, t_1590, t_1591);
not(t_1592, n41);
not(t_1593, g42);
and(c43, t_1592, t_1593);
not(t_1594, b42);
not(t_1595, j7);
and(d43, t_1594, t_1595);
not(t_1596, n39);
not(t_1597, c42);
and(e43, t_1596, t_1597);
not(t_1598, o41);
not(t_1599, h42);
and(f43, t_1598, t_1599);
not(t_1600, c42);
not(t_1601, z7);
and(g43, t_1600, t_1601);
not(t_1602, o39);
not(t_1603, d42);
and(h43, t_1602, t_1603);
not(t_1604, p41);
not(t_1605, i42);
and(i43, t_1604, t_1605);
not(t_1606, d42);
not(t_1607, p8);
and(j43, t_1606, t_1607);
not(t_1608, p39);
not(t_1609, e42);
and(k43, t_1608, t_1609);
not(t_1610, q41);
not(t_1611, j42);
and(l43, t_1610, t_1611);
not(t_1612, e42);
not(t_1613, f9);
and(m43, t_1612, t_1613);
not(t_1614, q39);
not(t_1615, f42);
and(n43, t_1614, t_1615);
not(t_1616, f42);
not(t_1617, v9);
and(o43, t_1616, t_1617);
not(t_1618, r39);
not(t_1619, g42);
and(p43, t_1618, t_1619);
not(t_1620, g42);
not(t_1621, l10);
and(q43, t_1620, t_1621);
not(t_1622, s39);
not(t_1623, h42);
and(r43, t_1622, t_1623);
not(t_1624, h42);
not(t_1625, b11);
and(s43, t_1624, t_1625);
not(t_1626, t39);
not(t_1627, i42);
and(t43, t_1626, t_1627);
not(t_1628, i42);
not(t_1629, r11);
and(u43, t_1628, t_1629);
not(t_1630, u39);
not(t_1631, j42);
and(v43, t_1630, t_1631);
not(t_1632, j42);
not(t_1633, h12);
and(w43, t_1632, t_1633);
not(t_1634, a3);
not(t_1635, k42);
and(x43, t_1634, t_1635);
not(t_1636, l42);
not(t_1637, s42);
and(y43, t_1636, t_1637);
not(t_1638, x39);
not(t_1639, u42);
and(z43, t_1638, t_1639);
not(t_1640, r41);
not(t_1641, u42);
and(a44, t_1640, t_1641);
not(t_1642, n42);
not(t_1643, o42);
and(b44, t_1642, t_1643);
not(t_1644, v41);
not(t_1645, p42);
and(c44, t_1644, t_1645);
not(t_1646, p42);
not(t_1647, w41);
and(d44, t_1646, t_1647);
not(t_1648, q42);
not(t_1649, y42);
and(e44, t_1648, t_1649);
not(t_1650, r42);
not(t_1651, a43);
and(f44, t_1650, t_1651);
not(t_1652, t42);
not(t_1653, d43);
and(g44, t_1652, t_1653);
not(t_1654, u42);
not(t_1655, g4);
and(h44, t_1654, t_1655);
not(t_1656, v42);
not(t_1657, g43);
and(i44, t_1656, t_1657);
not(t_1658, m42);
not(t_1659, w4);
and(j44, t_1658, t_1659);
not(t_1660, w42);
not(t_1661, j43);
and(k44, t_1660, t_1661);
not(t_1662, x42);
not(t_1663, m43);
and(l44, t_1662, t_1663);
not(t_1664, z42);
not(t_1665, o43);
and(m44, t_1664, t_1665);
not(t_1666, c43);
not(t_1667, q43);
and(n44, t_1666, t_1667);
not(t_1668, f43);
not(t_1669, s43);
and(o44, t_1668, t_1669);
not(t_1670, i43);
not(t_1671, u43);
and(p44, t_1670, t_1671);
not(t_1672, a3);
not(t_1673, x43);
and(q44, t_1672, t_1673);
not(t_1674, x43);
not(t_1675, k42);
and(r44, t_1674, t_1675);
not(t_1676, y43);
not(t_1677, z43);
and(s44, t_1676, t_1677);
not(t_1678, a44);
not(t_1679, h44);
and(t44, t_1678, t_1679);
not(t_1680, b41);
not(t_1681, j44);
and(u44, t_1680, t_1681);
not(t_1682, m42);
not(t_1683, j44);
and(v44, t_1682, t_1683);
not(t_1684, c44);
not(t_1685, d44);
and(w44, t_1684, t_1685);
not(t_1686, q42);
not(t_1687, e44);
and(x44, t_1686, t_1687);
not(t_1688, j44);
not(t_1689, w4);
and(y44, t_1688, t_1689);
not(t_1690, b44);
not(t_1691, m5);
and(z44, t_1690, t_1691);
not(t_1692, e44);
not(t_1693, y42);
and(a45, t_1692, t_1693);
not(t_1694, f44);
not(t_1695, b43);
and(b45, t_1694, t_1695);
not(t_1696, g44);
not(t_1697, e43);
and(c45, t_1696, t_1697);
not(t_1698, i44);
not(t_1699, h43);
and(d45, t_1698, t_1699);
not(t_1700, k44);
not(t_1701, k43);
and(e45, t_1700, t_1701);
not(t_1702, l44);
not(t_1703, n43);
and(f45, t_1702, t_1703);
not(t_1704, m44);
not(t_1705, p43);
and(g45, t_1704, t_1705);
not(t_1706, n44);
not(t_1707, r43);
and(h45, t_1706, t_1707);
not(t_1708, o44);
not(t_1709, t43);
and(i45, t_1708, t_1709);
not(t_1710, p44);
not(t_1711, v43);
and(j45, t_1710, t_1711);
not(t_1712, q44);
not(t_1713, r44);
and(k45, t_1712, t_1713);
not(t_1714, y43);
not(t_1715, s44);
and(l45, t_1714, t_1715);
not(t_1716, s44);
not(t_1717, z43);
and(m45, t_1716, t_1717);
not(t_1718, t44);
not(t_1719, u44);
and(n45, t_1718, t_1719);
not(t_1720, v44);
not(t_1721, y44);
and(o45, t_1720, t_1721);
not(t_1722, u41);
not(t_1723, z44);
and(p45, t_1722, t_1723);
not(t_1724, b44);
not(t_1725, z44);
and(q45, t_1724, t_1725);
not(t_1726, x44);
not(t_1727, a45);
and(r45, t_1726, t_1727);
not(t_1728, f44);
not(t_1729, b45);
and(s45, t_1728, t_1729);
not(t_1730, g44);
not(t_1731, c45);
and(t45, t_1730, t_1731);
not(t_1732, i44);
not(t_1733, d45);
and(u45, t_1732, t_1733);
not(t_1734, k44);
not(t_1735, e45);
and(v45, t_1734, t_1735);
not(t_1736, z44);
not(t_1737, m5);
and(w45, t_1736, t_1737);
not(t_1738, l44);
not(t_1739, f45);
and(x45, t_1738, t_1739);
not(t_1740, w44);
not(t_1741, c6);
and(y45, t_1740, t_1741);
not(t_1742, m44);
not(t_1743, g45);
and(z45, t_1742, t_1743);
not(t_1744, b45);
not(t_1745, b43);
and(a46, t_1744, t_1745);
not(t_1746, n44);
not(t_1747, h45);
and(b46, t_1746, t_1747);
not(t_1748, c45);
not(t_1749, e43);
and(c46, t_1748, t_1749);
not(t_1750, o44);
not(t_1751, i45);
and(d46, t_1750, t_1751);
not(t_1752, d45);
not(t_1753, h43);
and(e46, t_1752, t_1753);
not(t_1754, p44);
not(t_1755, j45);
and(f46, t_1754, t_1755);
not(t_1756, e45);
not(t_1757, k43);
and(g46, t_1756, t_1757);
not(t_1758, f45);
not(t_1759, n43);
and(h46, t_1758, t_1759);
not(t_1760, g45);
not(t_1761, p43);
and(i46, t_1760, t_1761);
not(t_1762, h45);
not(t_1763, r43);
and(j46, t_1762, t_1763);
not(t_1764, i45);
not(t_1765, t43);
and(k46, t_1764, t_1765);
not(t_1766, j45);
not(t_1767, v43);
and(l46, t_1766, t_1767);
not(t_1768, l45);
not(t_1769, m45);
and(m46, t_1768, t_1769);
not(t_1770, t44);
not(t_1771, n45);
and(n46, t_1770, t_1771);
not(t_1772, n45);
not(t_1773, u44);
and(o46, t_1772, t_1773);
not(t_1774, o45);
not(t_1775, p45);
and(p46, t_1774, t_1775);
not(t_1776, q45);
not(t_1777, w45);
and(q46, t_1776, t_1777);
not(t_1778, p42);
not(t_1779, y45);
and(r46, t_1778, t_1779);
not(t_1780, w44);
not(t_1781, y45);
and(s46, t_1780, t_1781);
not(t_1782, s45);
not(t_1783, a46);
and(t46, t_1782, t_1783);
not(t_1784, k45);
not(t_1785, p3);
and(u46, t_1784, t_1785);
not(t_1786, t45);
not(t_1787, c46);
and(v46, t_1786, t_1787);
not(t_1788, u45);
not(t_1789, e46);
and(w46, t_1788, t_1789);
not(t_1790, v45);
not(t_1791, g46);
and(x46, t_1790, t_1791);
not(t_1792, x45);
not(t_1793, h46);
and(y46, t_1792, t_1793);
not(t_1794, y45);
not(t_1795, c6);
and(z46, t_1794, t_1795);
not(t_1796, z45);
not(t_1797, i46);
and(a47, t_1796, t_1797);
not(t_1798, r45);
not(t_1799, s6);
and(b47, t_1798, t_1799);
not(t_1800, b46);
not(t_1801, j46);
and(c47, t_1800, t_1801);
not(t_1802, d46);
not(t_1803, k46);
and(d47, t_1802, t_1803);
not(t_1804, f46);
not(t_1805, l46);
and(e47, t_1804, t_1805);
not(t_1806, x43);
not(t_1807, u46);
and(f47, t_1806, t_1807);
not(t_1808, k45);
not(t_1809, u46);
and(g47, t_1808, t_1809);
not(t_1810, n46);
not(t_1811, o46);
and(h47, t_1810, t_1811);
not(t_1812, o45);
not(t_1813, p46);
and(i47, t_1812, t_1813);
not(t_1814, p46);
not(t_1815, p45);
and(j47, t_1814, t_1815);
not(t_1816, q46);
not(t_1817, r46);
and(k47, t_1816, t_1817);
not(t_1818, s46);
not(t_1819, z46);
and(l47, t_1818, t_1819);
not(t_1820, e44);
not(t_1821, b47);
and(m47, t_1820, t_1821);
not(t_1822, r45);
not(t_1823, b47);
and(n47, t_1822, t_1823);
not(t_1824, u46);
not(t_1825, p3);
and(o47, t_1824, t_1825);
not(t_1826, m46);
not(t_1827, f4);
and(p47, t_1826, t_1827);
not(t_1828, b47);
not(t_1829, s6);
and(q47, t_1828, t_1829);
not(t_1830, t46);
not(t_1831, i7);
and(r47, t_1830, t_1831);
not(t_1832, v46);
not(t_1833, y7);
and(s47, t_1832, t_1833);
not(t_1834, w46);
not(t_1835, o8);
and(t47, t_1834, t_1835);
not(t_1836, x46);
not(t_1837, e9);
and(u47, t_1836, t_1837);
not(t_1838, y46);
not(t_1839, u9);
and(v47, t_1838, t_1839);
not(t_1840, a47);
not(t_1841, k10);
and(w47, t_1840, t_1841);
not(t_1842, c47);
not(t_1843, a11);
and(x47, t_1842, t_1843);
not(t_1844, d47);
not(t_1845, q11);
and(y47, t_1844, t_1845);
not(t_1846, e47);
not(t_1847, g12);
and(z47, t_1846, t_1847);
not(t_1848, z2);
not(t_1849, f47);
and(a48, t_1848, t_1849);
not(t_1850, g47);
not(t_1851, o47);
and(b48, t_1850, t_1851);
not(t_1852, s44);
not(t_1853, p47);
and(c48, t_1852, t_1853);
not(t_1854, m46);
not(t_1855, p47);
and(d48, t_1854, t_1855);
not(t_1856, i47);
not(t_1857, j47);
and(e48, t_1856, t_1857);
not(t_1858, q46);
not(t_1859, k47);
and(f48, t_1858, t_1859);
not(t_1860, k47);
not(t_1861, r46);
and(g48, t_1860, t_1861);
not(t_1862, l47);
not(t_1863, m47);
and(h48, t_1862, t_1863);
not(t_1864, n47);
not(t_1865, q47);
and(i48, t_1864, t_1865);
not(t_1866, t46);
not(t_1867, r47);
and(j48, t_1866, t_1867);
not(t_1868, v46);
not(t_1869, s47);
and(k48, t_1868, t_1869);
not(t_1870, p47);
not(t_1871, f4);
and(l48, t_1870, t_1871);
not(t_1872, w46);
not(t_1873, t47);
and(m48, t_1872, t_1873);
not(t_1874, h47);
not(t_1875, v4);
and(n48, t_1874, t_1875);
not(t_1876, x46);
not(t_1877, u47);
and(o48, t_1876, t_1877);
not(t_1878, y46);
not(t_1879, v47);
and(p48, t_1878, t_1879);
not(t_1880, a47);
not(t_1881, w47);
and(q48, t_1880, t_1881);
not(t_1882, b45);
not(t_1883, r47);
and(r48, t_1882, t_1883);
not(t_1884, c47);
not(t_1885, x47);
and(s48, t_1884, t_1885);
not(t_1886, r47);
not(t_1887, i7);
and(t48, t_1886, t_1887);
not(t_1888, c45);
not(t_1889, s47);
and(u48, t_1888, t_1889);
not(t_1890, d47);
not(t_1891, y47);
and(v48, t_1890, t_1891);
not(t_1892, s47);
not(t_1893, y7);
and(w48, t_1892, t_1893);
not(t_1894, d45);
not(t_1895, t47);
and(x48, t_1894, t_1895);
not(t_1896, e47);
not(t_1897, z47);
and(y48, t_1896, t_1897);
not(t_1898, t47);
not(t_1899, o8);
and(z48, t_1898, t_1899);
not(t_1900, e45);
not(t_1901, u47);
and(a49, t_1900, t_1901);
not(t_1902, u47);
not(t_1903, e9);
and(b49, t_1902, t_1903);
not(t_1904, f45);
not(t_1905, v47);
and(c49, t_1904, t_1905);
not(t_1906, v47);
not(t_1907, u9);
and(d49, t_1906, t_1907);
not(t_1908, g45);
not(t_1909, w47);
and(e49, t_1908, t_1909);
not(t_1910, w47);
not(t_1911, k10);
and(f49, t_1910, t_1911);
not(t_1912, h45);
not(t_1913, x47);
and(g49, t_1912, t_1913);
not(t_1914, x47);
not(t_1915, a11);
and(h49, t_1914, t_1915);
not(t_1916, i45);
not(t_1917, y47);
and(i49, t_1916, t_1917);
not(t_1918, y47);
not(t_1919, q11);
and(j49, t_1918, t_1919);
not(t_1920, j45);
not(t_1921, z47);
and(k49, t_1920, t_1921);
not(t_1922, z47);
not(t_1923, g12);
and(l49, t_1922, t_1923);
not(t_1924, z2);
not(t_1925, a48);
and(m49, t_1924, t_1925);
not(t_1926, a48);
not(t_1927, f47);
and(n49, t_1926, t_1927);
not(t_1928, b48);
not(t_1929, c48);
and(o49, t_1928, t_1929);
not(t_1930, d48);
not(t_1931, l48);
and(p49, t_1930, t_1931);
not(t_1932, n45);
not(t_1933, n48);
and(q49, t_1932, t_1933);
not(t_1934, h47);
not(t_1935, n48);
and(r49, t_1934, t_1935);
not(t_1936, f48);
not(t_1937, g48);
and(s49, t_1936, t_1937);
not(t_1938, l47);
not(t_1939, h48);
and(t49, t_1938, t_1939);
not(t_1940, h48);
not(t_1941, m47);
and(u49, t_1940, t_1941);
not(t_1942, i48);
not(t_1943, r48);
and(v49, t_1942, t_1943);
not(t_1944, j48);
not(t_1945, t48);
and(w49, t_1944, t_1945);
not(t_1946, k48);
not(t_1947, w48);
and(x49, t_1946, t_1947);
not(t_1948, m48);
not(t_1949, z48);
and(y49, t_1948, t_1949);
not(t_1950, n48);
not(t_1951, v4);
and(z49, t_1950, t_1951);
not(t_1952, o48);
not(t_1953, b49);
and(a50, t_1952, t_1953);
not(t_1954, e48);
not(t_1955, l5);
and(b50, t_1954, t_1955);
not(t_1956, p48);
not(t_1957, d49);
and(c50, t_1956, t_1957);
not(t_1958, q48);
not(t_1959, f49);
and(d50, t_1958, t_1959);
not(t_1960, s48);
not(t_1961, h49);
and(e50, t_1960, t_1961);
not(t_1962, v48);
not(t_1963, j49);
and(f50, t_1962, t_1963);
not(t_1964, m49);
not(t_1965, n49);
and(g50, t_1964, t_1965);
not(t_1966, b48);
not(t_1967, o49);
and(h50, t_1966, t_1967);
not(t_1968, o49);
not(t_1969, c48);
and(i50, t_1968, t_1969);
not(t_1970, p49);
not(t_1971, q49);
and(j50, t_1970, t_1971);
not(t_1972, r49);
not(t_1973, z49);
and(k50, t_1972, t_1973);
not(t_1974, p46);
not(t_1975, b50);
and(l50, t_1974, t_1975);
not(t_1976, e48);
not(t_1977, b50);
and(m50, t_1976, t_1977);
not(t_1978, t49);
not(t_1979, u49);
and(n50, t_1978, t_1979);
not(t_1980, i48);
not(t_1981, v49);
and(o50, t_1980, t_1981);
not(t_1982, b50);
not(t_1983, l5);
and(p50, t_1982, t_1983);
not(t_1984, s49);
not(t_1985, b6);
and(q50, t_1984, t_1985);
not(t_1986, v49);
not(t_1987, r48);
and(r50, t_1986, t_1987);
not(t_1988, w49);
not(t_1989, u48);
and(s50, t_1988, t_1989);
not(t_1990, x49);
not(t_1991, x48);
and(t50, t_1990, t_1991);
not(t_1992, y49);
not(t_1993, a49);
and(u50, t_1992, t_1993);
not(t_1994, a50);
not(t_1995, c49);
and(v50, t_1994, t_1995);
not(t_1996, c50);
not(t_1997, e49);
and(w50, t_1996, t_1997);
not(t_1998, d50);
not(t_1999, g49);
and(x50, t_1998, t_1999);
not(t_2000, e50);
not(t_2001, i49);
and(y50, t_2000, t_2001);
not(t_2002, f50);
not(t_2003, k49);
and(z50, t_2002, t_2003);
not(t_2004, h50);
not(t_2005, i50);
and(a51, t_2004, t_2005);
not(t_2006, p49);
not(t_2007, j50);
and(b51, t_2006, t_2007);
not(t_2008, j50);
not(t_2009, q49);
and(c51, t_2008, t_2009);
not(t_2010, k50);
not(t_2011, l50);
and(d51, t_2010, t_2011);
not(t_2012, m50);
not(t_2013, p50);
and(e51, t_2012, t_2013);
not(t_2014, k47);
not(t_2015, q50);
and(f51, t_2014, t_2015);
not(t_2016, s49);
not(t_2017, q50);
and(g51, t_2016, t_2017);
not(t_2018, o50);
not(t_2019, r50);
and(h51, t_2018, t_2019);
not(t_2020, w49);
not(t_2021, s50);
and(i51, t_2020, t_2021);
not(t_2022, g50);
not(t_2023, o3);
and(j51, t_2022, t_2023);
not(t_2024, x49);
not(t_2025, t50);
and(k51, t_2024, t_2025);
not(t_2026, y49);
not(t_2027, u50);
and(l51, t_2026, t_2027);
not(t_2028, a50);
not(t_2029, v50);
and(m51, t_2028, t_2029);
not(t_2030, c50);
not(t_2031, w50);
and(n51, t_2030, t_2031);
not(t_2032, q50);
not(t_2033, b6);
and(o51, t_2032, t_2033);
not(t_2034, d50);
not(t_2035, x50);
and(p51, t_2034, t_2035);
not(t_2036, n50);
not(t_2037, r6);
and(q51, t_2036, t_2037);
not(t_2038, e50);
not(t_2039, y50);
and(r51, t_2038, t_2039);
not(t_2040, s50);
not(t_2041, u48);
and(s51, t_2040, t_2041);
not(t_2042, f50);
not(t_2043, z50);
and(t51, t_2042, t_2043);
not(t_2044, t50);
not(t_2045, x48);
and(u51, t_2044, t_2045);
not(t_2046, u50);
not(t_2047, a49);
and(v51, t_2046, t_2047);
not(t_2048, v50);
not(t_2049, c49);
and(w51, t_2048, t_2049);
not(t_2050, w50);
not(t_2051, e49);
and(x51, t_2050, t_2051);
not(t_2052, x50);
not(t_2053, g49);
and(y51, t_2052, t_2053);
not(t_2054, y50);
not(t_2055, i49);
and(z51, t_2054, t_2055);
not(t_2056, z50);
not(t_2057, k49);
and(a52, t_2056, t_2057);
not(t_2058, a48);
not(t_2059, j51);
and(b52, t_2058, t_2059);
not(t_2060, g50);
not(t_2061, j51);
and(c52, t_2060, t_2061);
not(t_2062, b51);
not(t_2063, c51);
and(d52, t_2062, t_2063);
not(t_2064, k50);
not(t_2065, d51);
and(e52, t_2064, t_2065);
not(t_2066, d51);
not(t_2067, l50);
and(f52, t_2066, t_2067);
not(t_2068, e51);
not(t_2069, f51);
and(g52, t_2068, t_2069);
not(t_2070, g51);
not(t_2071, o51);
and(h52, t_2070, t_2071);
not(t_2072, h48);
not(t_2073, q51);
and(i52, t_2072, t_2073);
not(t_2074, n50);
not(t_2075, q51);
and(j52, t_2074, t_2075);
not(t_2076, i51);
not(t_2077, s51);
and(k52, t_2076, t_2077);
not(t_2078, j51);
not(t_2079, o3);
and(l52, t_2078, t_2079);
not(t_2080, k51);
not(t_2081, u51);
and(m52, t_2080, t_2081);
not(t_2082, a51);
not(t_2083, e4);
and(n52, t_2082, t_2083);
not(t_2084, l51);
not(t_2085, v51);
and(o52, t_2084, t_2085);
not(t_2086, m51);
not(t_2087, w51);
and(p52, t_2086, t_2087);
not(t_2088, n51);
not(t_2089, x51);
and(q52, t_2088, t_2089);
not(t_2090, p51);
not(t_2091, y51);
and(r52, t_2090, t_2091);
not(t_2092, q51);
not(t_2093, r6);
and(s52, t_2092, t_2093);
not(t_2094, r51);
not(t_2095, z51);
and(t52, t_2094, t_2095);
not(t_2096, h51);
not(t_2097, h7);
and(u52, t_2096, t_2097);
not(t_2098, t51);
not(t_2099, a52);
and(v52, t_2098, t_2099);
not(t_2100, y2);
not(t_2101, b52);
and(w52, t_2100, t_2101);
not(t_2102, c52);
not(t_2103, l52);
and(x52, t_2102, t_2103);
not(t_2104, o49);
not(t_2105, n52);
and(y52, t_2104, t_2105);
not(t_2106, a51);
not(t_2107, n52);
and(z52, t_2106, t_2107);
not(t_2108, e52);
not(t_2109, f52);
and(a53, t_2108, t_2109);
not(t_2110, e51);
not(t_2111, g52);
and(b53, t_2110, t_2111);
not(t_2112, g52);
not(t_2113, f51);
and(c53, t_2112, t_2113);
not(t_2114, h52);
not(t_2115, i52);
and(d53, t_2114, t_2115);
not(t_2116, j52);
not(t_2117, s52);
and(e53, t_2116, t_2117);
not(t_2118, v49);
not(t_2119, u52);
and(f53, t_2118, t_2119);
not(t_2120, h51);
not(t_2121, u52);
and(g53, t_2120, t_2121);
not(t_2122, n52);
not(t_2123, e4);
and(h53, t_2122, t_2123);
not(t_2124, d52);
not(t_2125, u4);
and(i53, t_2124, t_2125);
not(t_2126, u52);
not(t_2127, h7);
and(j53, t_2126, t_2127);
not(t_2128, k52);
not(t_2129, x7);
and(k53, t_2128, t_2129);
not(t_2130, m52);
not(t_2131, n8);
and(l53, t_2130, t_2131);
not(t_2132, o52);
not(t_2133, d9);
and(m53, t_2132, t_2133);
not(t_2134, p52);
not(t_2135, t9);
and(n53, t_2134, t_2135);
not(t_2136, q52);
not(t_2137, j10);
and(o53, t_2136, t_2137);
not(t_2138, r52);
not(t_2139, z10);
and(p53, t_2138, t_2139);
not(t_2140, t52);
not(t_2141, p11);
and(q53, t_2140, t_2141);
not(t_2142, v52);
not(t_2143, f12);
and(r53, t_2142, t_2143);
not(t_2144, y2);
not(t_2145, w52);
and(s53, t_2144, t_2145);
not(t_2146, w52);
not(t_2147, b52);
and(t53, t_2146, t_2147);
not(t_2148, x52);
not(t_2149, y52);
and(u53, t_2148, t_2149);
not(t_2150, z52);
not(t_2151, h53);
and(v53, t_2150, t_2151);
not(t_2152, j50);
not(t_2153, i53);
and(w53, t_2152, t_2153);
not(t_2154, d52);
not(t_2155, i53);
and(x53, t_2154, t_2155);
not(t_2156, b53);
not(t_2157, c53);
and(y53, t_2156, t_2157);
not(t_2158, h52);
not(t_2159, d53);
and(z53, t_2158, t_2159);
not(t_2160, d53);
not(t_2161, i52);
and(a54, t_2160, t_2161);
not(t_2162, e53);
not(t_2163, f53);
and(b54, t_2162, t_2163);
not(t_2164, g53);
not(t_2165, j53);
and(c54, t_2164, t_2165);
not(t_2166, k52);
not(t_2167, k53);
and(d54, t_2166, t_2167);
not(t_2168, m52);
not(t_2169, l53);
and(e54, t_2168, t_2169);
not(t_2170, o52);
not(t_2171, m53);
and(f54, t_2170, t_2171);
not(t_2172, i53);
not(t_2173, u4);
and(g54, t_2172, t_2173);
not(t_2174, p52);
not(t_2175, n53);
and(h54, t_2174, t_2175);
not(t_2176, a53);
not(t_2177, k5);
and(i54, t_2176, t_2177);
not(t_2178, q52);
not(t_2179, o53);
and(j54, t_2178, t_2179);
not(t_2180, r52);
not(t_2181, p53);
and(k54, t_2180, t_2181);
not(t_2182, t52);
not(t_2183, q53);
and(l54, t_2182, t_2183);
not(t_2184, s50);
not(t_2185, k53);
and(m54, t_2184, t_2185);
not(t_2186, v52);
not(t_2187, r53);
and(n54, t_2186, t_2187);
not(t_2188, k53);
not(t_2189, x7);
and(o54, t_2188, t_2189);
not(t_2190, t50);
not(t_2191, l53);
and(p54, t_2190, t_2191);
not(t_2192, l53);
not(t_2193, n8);
and(q54, t_2192, t_2193);
not(t_2194, u50);
not(t_2195, m53);
and(r54, t_2194, t_2195);
not(t_2196, m53);
not(t_2197, d9);
and(s54, t_2196, t_2197);
not(t_2198, v50);
not(t_2199, n53);
and(t54, t_2198, t_2199);
not(t_2200, n53);
not(t_2201, t9);
and(u54, t_2200, t_2201);
not(t_2202, w50);
not(t_2203, o53);
and(v54, t_2202, t_2203);
not(t_2204, o53);
not(t_2205, j10);
and(w54, t_2204, t_2205);
not(t_2206, x50);
not(t_2207, p53);
and(x54, t_2206, t_2207);
not(t_2208, p53);
not(t_2209, z10);
and(y54, t_2208, t_2209);
not(t_2210, y50);
not(t_2211, q53);
and(z54, t_2210, t_2211);
not(t_2212, q53);
not(t_2213, p11);
and(a55, t_2212, t_2213);
not(t_2214, z50);
not(t_2215, r53);
and(b55, t_2214, t_2215);
not(t_2216, r53);
not(t_2217, f12);
and(c55, t_2216, t_2217);
not(t_2218, s53);
not(t_2219, t53);
and(d55, t_2218, t_2219);
not(t_2220, x52);
not(t_2221, u53);
and(e55, t_2220, t_2221);
not(t_2222, u53);
not(t_2223, y52);
and(f55, t_2222, t_2223);
not(t_2224, v53);
not(t_2225, w53);
and(g55, t_2224, t_2225);
not(t_2226, x53);
not(t_2227, g54);
and(h55, t_2226, t_2227);
not(t_2228, d51);
not(t_2229, i54);
and(i55, t_2228, t_2229);
not(t_2230, a53);
not(t_2231, i54);
and(j55, t_2230, t_2231);
not(t_2232, z53);
not(t_2233, a54);
and(k55, t_2232, t_2233);
not(t_2234, e53);
not(t_2235, b54);
and(l55, t_2234, t_2235);
not(t_2236, b54);
not(t_2237, f53);
and(m55, t_2236, t_2237);
not(t_2238, c54);
not(t_2239, m54);
and(n55, t_2238, t_2239);
not(t_2240, d54);
not(t_2241, o54);
and(o55, t_2240, t_2241);
not(t_2242, e54);
not(t_2243, q54);
and(p55, t_2242, t_2243);
not(t_2244, f54);
not(t_2245, s54);
and(q55, t_2244, t_2245);
not(t_2246, h54);
not(t_2247, u54);
and(r55, t_2246, t_2247);
not(t_2248, i54);
not(t_2249, k5);
and(s55, t_2248, t_2249);
not(t_2250, j54);
not(t_2251, w54);
and(t55, t_2250, t_2251);
not(t_2252, y53);
not(t_2253, a6);
and(u55, t_2252, t_2253);
not(t_2254, k54);
not(t_2255, y54);
and(v55, t_2254, t_2255);
not(t_2256, l54);
not(t_2257, a55);
and(w55, t_2256, t_2257);
not(t_2258, e55);
not(t_2259, f55);
and(x55, t_2258, t_2259);
not(t_2260, v53);
not(t_2261, g55);
and(y55, t_2260, t_2261);
not(t_2262, g55);
not(t_2263, w53);
and(z55, t_2262, t_2263);
not(t_2264, h55);
not(t_2265, i55);
and(a56, t_2264, t_2265);
not(t_2266, j55);
not(t_2267, s55);
and(b56, t_2266, t_2267);
not(t_2268, g52);
not(t_2269, u55);
and(c56, t_2268, t_2269);
not(t_2270, y53);
not(t_2271, u55);
and(d56, t_2270, t_2271);
not(t_2272, l55);
not(t_2273, m55);
and(e56, t_2272, t_2273);
not(t_2274, c54);
not(t_2275, n55);
and(f56, t_2274, t_2275);
not(t_2276, d55);
not(t_2277, n3);
and(g56, t_2276, t_2277);
not(t_2278, u55);
not(t_2279, a6);
and(h56, t_2278, t_2279);
not(t_2280, k55);
not(t_2281, q6);
and(i56, t_2280, t_2281);
not(t_2282, n55);
not(t_2283, m54);
and(j56, t_2282, t_2283);
not(t_2284, o55);
not(t_2285, p54);
and(k56, t_2284, t_2285);
not(t_2286, p55);
not(t_2287, r54);
and(l56, t_2286, t_2287);
not(t_2288, q55);
not(t_2289, t54);
and(m56, t_2288, t_2289);
not(t_2290, r55);
not(t_2291, v54);
and(n56, t_2290, t_2291);
not(t_2292, t55);
not(t_2293, x54);
and(o56, t_2292, t_2293);
not(t_2294, v55);
not(t_2295, z54);
and(p56, t_2294, t_2295);
not(t_2296, w55);
not(t_2297, b55);
and(q56, t_2296, t_2297);
not(t_2298, w52);
not(t_2299, g56);
and(r56, t_2298, t_2299);
not(t_2300, d55);
not(t_2301, g56);
and(s56, t_2300, t_2301);
not(t_2302, y55);
not(t_2303, z55);
and(t56, t_2302, t_2303);
not(t_2304, h55);
not(t_2305, a56);
and(u56, t_2304, t_2305);
not(t_2306, a56);
not(t_2307, i55);
and(v56, t_2306, t_2307);
not(t_2308, b56);
not(t_2309, c56);
and(w56, t_2308, t_2309);
not(t_2310, d56);
not(t_2311, h56);
and(x56, t_2310, t_2311);
not(t_2312, d53);
not(t_2313, i56);
and(y56, t_2312, t_2313);
not(t_2314, k55);
not(t_2315, i56);
and(z56, t_2314, t_2315);
not(t_2316, f56);
not(t_2317, j56);
and(a57, t_2316, t_2317);
not(t_2318, o55);
not(t_2319, k56);
and(b57, t_2318, t_2319);
not(t_2320, g56);
not(t_2321, n3);
and(c57, t_2320, t_2321);
not(t_2322, p55);
not(t_2323, l56);
and(d57, t_2322, t_2323);
not(t_2324, x55);
not(t_2325, d4);
and(e57, t_2324, t_2325);
not(t_2326, q55);
not(t_2327, m56);
and(f57, t_2326, t_2327);
not(t_2328, r55);
not(t_2329, n56);
and(g57, t_2328, t_2329);
not(t_2330, t55);
not(t_2331, o56);
and(h57, t_2330, t_2331);
not(t_2332, v55);
not(t_2333, p56);
and(i57, t_2332, t_2333);
not(t_2334, i56);
not(t_2335, q6);
and(j57, t_2334, t_2335);
not(t_2336, w55);
not(t_2337, q56);
and(k57, t_2336, t_2337);
not(t_2338, e56);
not(t_2339, g7);
and(l57, t_2338, t_2339);
not(t_2340, k56);
not(t_2341, p54);
and(m57, t_2340, t_2341);
not(t_2342, l56);
not(t_2343, r54);
and(n57, t_2342, t_2343);
not(t_2344, m56);
not(t_2345, t54);
and(o57, t_2344, t_2345);
not(t_2346, n56);
not(t_2347, v54);
and(p57, t_2346, t_2347);
not(t_2348, o56);
not(t_2349, x54);
and(q57, t_2348, t_2349);
not(t_2350, p56);
not(t_2351, z54);
and(r57, t_2350, t_2351);
not(t_2352, q56);
not(t_2353, b55);
and(s57, t_2352, t_2353);
not(t_2354, x2);
not(t_2355, r56);
and(t57, t_2354, t_2355);
not(t_2356, s56);
not(t_2357, c57);
and(u57, t_2356, t_2357);
not(t_2358, u53);
not(t_2359, e57);
and(v57, t_2358, t_2359);
not(t_2360, x55);
not(t_2361, e57);
and(w57, t_2360, t_2361);
not(t_2362, u56);
not(t_2363, v56);
and(x57, t_2362, t_2363);
not(t_2364, b56);
not(t_2365, w56);
and(y57, t_2364, t_2365);
not(t_2366, w56);
not(t_2367, c56);
and(z57, t_2366, t_2367);
not(t_2368, x56);
not(t_2369, y56);
and(a58, t_2368, t_2369);
not(t_2370, z56);
not(t_2371, j57);
and(b58, t_2370, t_2371);
not(t_2372, b54);
not(t_2373, l57);
and(c58, t_2372, t_2373);
not(t_2374, e56);
not(t_2375, l57);
and(d58, t_2374, t_2375);
not(t_2376, b57);
not(t_2377, m57);
and(e58, t_2376, t_2377);
not(t_2378, d57);
not(t_2379, n57);
and(f58, t_2378, t_2379);
not(t_2380, e57);
not(t_2381, d4);
and(g58, t_2380, t_2381);
not(t_2382, f57);
not(t_2383, o57);
and(h58, t_2382, t_2383);
not(t_2384, t56);
not(t_2385, t4);
and(i58, t_2384, t_2385);
not(t_2386, g57);
not(t_2387, p57);
and(j58, t_2386, t_2387);
not(t_2388, h57);
not(t_2389, q57);
and(k58, t_2388, t_2389);
not(t_2390, i57);
not(t_2391, r57);
and(l58, t_2390, t_2391);
not(t_2392, k57);
not(t_2393, s57);
and(m58, t_2392, t_2393);
not(t_2394, l57);
not(t_2395, g7);
and(n58, t_2394, t_2395);
not(t_2396, a57);
not(t_2397, w7);
and(o58, t_2396, t_2397);
not(t_2398, x2);
not(t_2399, t57);
and(p58, t_2398, t_2399);
not(t_2400, t57);
not(t_2401, r56);
and(q58, t_2400, t_2401);
not(t_2402, u57);
not(t_2403, v57);
and(r58, t_2402, t_2403);
not(t_2404, w57);
not(t_2405, g58);
and(s58, t_2404, t_2405);
not(t_2406, g55);
not(t_2407, i58);
and(t58, t_2406, t_2407);
not(t_2408, t56);
not(t_2409, i58);
and(u58, t_2408, t_2409);
not(t_2410, y57);
not(t_2411, z57);
and(v58, t_2410, t_2411);
not(t_2412, x56);
not(t_2413, a58);
and(w58, t_2412, t_2413);
not(t_2414, a58);
not(t_2415, y56);
and(x58, t_2414, t_2415);
not(t_2416, b58);
not(t_2417, c58);
and(y58, t_2416, t_2417);
not(t_2418, d58);
not(t_2419, n58);
and(z58, t_2418, t_2419);
not(t_2420, n55);
not(t_2421, o58);
and(a59, t_2420, t_2421);
not(t_2422, a57);
not(t_2423, o58);
and(b59, t_2422, t_2423);
not(t_2424, i58);
not(t_2425, t4);
and(c59, t_2424, t_2425);
not(t_2426, x57);
not(t_2427, j5);
and(d59, t_2426, t_2427);
not(t_2428, o58);
not(t_2429, w7);
and(e59, t_2428, t_2429);
not(t_2430, e58);
not(t_2431, m8);
and(f59, t_2430, t_2431);
not(t_2432, f58);
not(t_2433, c9);
and(g59, t_2432, t_2433);
not(t_2434, h58);
not(t_2435, s9);
and(h59, t_2434, t_2435);
not(t_2436, j58);
not(t_2437, i10);
and(i59, t_2436, t_2437);
not(t_2438, k58);
not(t_2439, y10);
and(j59, t_2438, t_2439);
not(t_2440, l58);
not(t_2441, o11);
and(k59, t_2440, t_2441);
not(t_2442, m58);
not(t_2443, e12);
and(l59, t_2442, t_2443);
not(t_2444, p58);
not(t_2445, q58);
and(m59, t_2444, t_2445);
not(t_2446, u57);
not(t_2447, r58);
and(n59, t_2446, t_2447);
not(t_2448, r58);
not(t_2449, v57);
and(o59, t_2448, t_2449);
not(t_2450, s58);
not(t_2451, t58);
and(p59, t_2450, t_2451);
not(t_2452, u58);
not(t_2453, c59);
and(q59, t_2452, t_2453);
not(t_2454, a56);
not(t_2455, d59);
and(r59, t_2454, t_2455);
not(t_2456, x57);
not(t_2457, d59);
and(s59, t_2456, t_2457);
not(t_2458, w58);
not(t_2459, x58);
and(t59, t_2458, t_2459);
not(t_2460, b58);
not(t_2461, y58);
and(u59, t_2460, t_2461);
not(t_2462, y58);
not(t_2463, c58);
and(v59, t_2462, t_2463);
not(t_2464, z58);
not(t_2465, a59);
and(w59, t_2464, t_2465);
not(t_2466, b59);
not(t_2467, e59);
and(x59, t_2466, t_2467);
not(t_2468, e58);
not(t_2469, f59);
and(y59, t_2468, t_2469);
not(t_2470, f58);
not(t_2471, g59);
and(z59, t_2470, t_2471);
not(t_2472, h58);
not(t_2473, h59);
and(a60, t_2472, t_2473);
not(t_2474, j58);
not(t_2475, i59);
and(b60, t_2474, t_2475);
not(t_2476, d59);
not(t_2477, j5);
and(c60, t_2476, t_2477);
not(t_2478, k58);
not(t_2479, j59);
and(d60, t_2478, t_2479);
not(t_2480, v58);
not(t_2481, z5);
and(e60, t_2480, t_2481);
not(t_2482, l58);
not(t_2483, k59);
and(f60, t_2482, t_2483);
not(t_2484, m58);
not(t_2485, l59);
and(g60, t_2484, t_2485);
not(t_2486, k56);
not(t_2487, f59);
and(h60, t_2486, t_2487);
not(t_2488, f59);
not(t_2489, m8);
and(i60, t_2488, t_2489);
not(t_2490, l56);
not(t_2491, g59);
and(j60, t_2490, t_2491);
not(t_2492, g59);
not(t_2493, c9);
and(k60, t_2492, t_2493);
not(t_2494, m56);
not(t_2495, h59);
and(l60, t_2494, t_2495);
not(t_2496, h59);
not(t_2497, s9);
and(m60, t_2496, t_2497);
not(t_2498, n56);
not(t_2499, i59);
and(n60, t_2498, t_2499);
not(t_2500, i59);
not(t_2501, i10);
and(o60, t_2500, t_2501);
not(t_2502, o56);
not(t_2503, j59);
and(p60, t_2502, t_2503);
not(t_2504, j59);
not(t_2505, y10);
and(q60, t_2504, t_2505);
not(t_2506, p56);
not(t_2507, k59);
and(r60, t_2506, t_2507);
not(t_2508, k59);
not(t_2509, o11);
and(s60, t_2508, t_2509);
not(t_2510, q56);
not(t_2511, l59);
and(t60, t_2510, t_2511);
not(t_2512, l59);
not(t_2513, e12);
and(u60, t_2512, t_2513);
not(t_2514, n59);
not(t_2515, o59);
and(v60, t_2514, t_2515);
not(t_2516, s58);
not(t_2517, p59);
and(w60, t_2516, t_2517);
not(t_2518, p59);
not(t_2519, t58);
and(x60, t_2518, t_2519);
not(t_2520, q59);
not(t_2521, r59);
and(y60, t_2520, t_2521);
not(t_2522, s59);
not(t_2523, c60);
and(z60, t_2522, t_2523);
not(t_2524, w56);
not(t_2525, e60);
and(a61, t_2524, t_2525);
not(t_2526, v58);
not(t_2527, e60);
and(b61, t_2526, t_2527);
not(t_2528, u59);
not(t_2529, v59);
and(c61, t_2528, t_2529);
not(t_2530, z58);
not(t_2531, w59);
and(d61, t_2530, t_2531);
not(t_2532, w59);
not(t_2533, a59);
and(e61, t_2532, t_2533);
not(t_2534, x59);
not(t_2535, h60);
and(f61, t_2534, t_2535);
not(t_2536, y59);
not(t_2537, i60);
and(g61, t_2536, t_2537);
not(t_2538, m59);
not(t_2539, m3);
and(h61, t_2538, t_2539);
not(t_2540, z59);
not(t_2541, k60);
and(i61, t_2540, t_2541);
not(t_2542, a60);
not(t_2543, m60);
and(j61, t_2542, t_2543);
not(t_2544, b60);
not(t_2545, o60);
and(k61, t_2544, t_2545);
not(t_2546, d60);
not(t_2547, q60);
and(l61, t_2546, t_2547);
not(t_2548, e60);
not(t_2549, z5);
and(m61, t_2548, t_2549);
not(t_2550, f60);
not(t_2551, s60);
and(n61, t_2550, t_2551);
not(t_2552, t59);
not(t_2553, p6);
and(o61, t_2552, t_2553);
not(t_2554, t57);
not(t_2555, h61);
and(p61, t_2554, t_2555);
not(t_2556, m59);
not(t_2557, h61);
and(q61, t_2556, t_2557);
not(t_2558, w60);
not(t_2559, x60);
and(r61, t_2558, t_2559);
not(t_2560, q59);
not(t_2561, y60);
and(s61, t_2560, t_2561);
not(t_2562, y60);
not(t_2563, r59);
and(t61, t_2562, t_2563);
not(t_2564, z60);
not(t_2565, a61);
and(u61, t_2564, t_2565);
not(t_2566, b61);
not(t_2567, m61);
and(v61, t_2566, t_2567);
not(t_2568, a58);
not(t_2569, o61);
and(w61, t_2568, t_2569);
not(t_2570, t59);
not(t_2571, o61);
and(x61, t_2570, t_2571);
not(t_2572, d61);
not(t_2573, e61);
and(y61, t_2572, t_2573);
not(t_2574, x59);
not(t_2575, f61);
and(z61, t_2574, t_2575);
not(t_2576, h61);
not(t_2577, m3);
and(a62, t_2576, t_2577);
not(t_2578, v60);
not(t_2579, c4);
and(b62, t_2578, t_2579);
not(t_2580, o61);
not(t_2581, p6);
and(c62, t_2580, t_2581);
not(t_2582, c61);
not(t_2583, f7);
and(d62, t_2582, t_2583);
not(t_2584, f61);
not(t_2585, h60);
and(e62, t_2584, t_2585);
not(t_2586, g61);
not(t_2587, j60);
and(f62, t_2586, t_2587);
not(t_2588, i61);
not(t_2589, l60);
and(g62, t_2588, t_2589);
not(t_2590, j61);
not(t_2591, n60);
and(h62, t_2590, t_2591);
not(t_2592, k61);
not(t_2593, p60);
and(i62, t_2592, t_2593);
not(t_2594, l61);
not(t_2595, r60);
and(j62, t_2594, t_2595);
not(t_2596, n61);
not(t_2597, t60);
and(k62, t_2596, t_2597);
not(t_2598, w2);
not(t_2599, p61);
and(l62, t_2598, t_2599);
not(t_2600, q61);
not(t_2601, a62);
and(m62, t_2600, t_2601);
not(t_2602, r58);
not(t_2603, b62);
and(n62, t_2602, t_2603);
not(t_2604, v60);
not(t_2605, b62);
and(o62, t_2604, t_2605);
not(t_2606, s61);
not(t_2607, t61);
and(p62, t_2606, t_2607);
not(t_2608, z60);
not(t_2609, u61);
and(q62, t_2608, t_2609);
not(t_2610, u61);
not(t_2611, a61);
and(r62, t_2610, t_2611);
not(t_2612, v61);
not(t_2613, w61);
and(s62, t_2612, t_2613);
not(t_2614, x61);
not(t_2615, c62);
and(t62, t_2614, t_2615);
not(t_2616, y58);
not(t_2617, d62);
and(u62, t_2616, t_2617);
not(t_2618, c61);
not(t_2619, d62);
and(v62, t_2618, t_2619);
not(t_2620, z61);
not(t_2621, e62);
and(w62, t_2620, t_2621);
not(t_2622, g61);
not(t_2623, f62);
and(x62, t_2622, t_2623);
not(t_2624, i61);
not(t_2625, g62);
and(y62, t_2624, t_2625);
not(t_2626, b62);
not(t_2627, c4);
and(z62, t_2626, t_2627);
not(t_2628, j61);
not(t_2629, h62);
and(a63, t_2628, t_2629);
not(t_2630, r61);
not(t_2631, s4);
and(b63, t_2630, t_2631);
not(t_2632, k61);
not(t_2633, i62);
and(c63, t_2632, t_2633);
not(t_2634, l61);
not(t_2635, j62);
and(d63, t_2634, t_2635);
not(t_2636, n61);
not(t_2637, k62);
and(e63, t_2636, t_2637);
not(t_2638, d62);
not(t_2639, f7);
and(f63, t_2638, t_2639);
not(t_2640, y61);
not(t_2641, v7);
and(g63, t_2640, t_2641);
not(t_2642, f62);
not(t_2643, j60);
and(h63, t_2642, t_2643);
not(t_2644, g62);
not(t_2645, l60);
and(i63, t_2644, t_2645);
not(t_2646, h62);
not(t_2647, n60);
and(j63, t_2646, t_2647);
not(t_2648, i62);
not(t_2649, p60);
and(k63, t_2648, t_2649);
not(t_2650, j62);
not(t_2651, r60);
and(l63, t_2650, t_2651);
not(t_2652, k62);
not(t_2653, t60);
and(m63, t_2652, t_2653);
not(t_2654, w2);
not(t_2655, l62);
and(n63, t_2654, t_2655);
not(t_2656, l62);
not(t_2657, p61);
and(o63, t_2656, t_2657);
not(t_2658, m62);
not(t_2659, n62);
and(p63, t_2658, t_2659);
not(t_2660, o62);
not(t_2661, z62);
and(q63, t_2660, t_2661);
not(t_2662, p59);
not(t_2663, b63);
and(r63, t_2662, t_2663);
not(t_2664, r61);
not(t_2665, b63);
and(s63, t_2664, t_2665);
not(t_2666, q62);
not(t_2667, r62);
and(t63, t_2666, t_2667);
not(t_2668, v61);
not(t_2669, s62);
and(u63, t_2668, t_2669);
not(t_2670, s62);
not(t_2671, w61);
and(v63, t_2670, t_2671);
not(t_2672, t62);
not(t_2673, u62);
and(w63, t_2672, t_2673);
not(t_2674, v62);
not(t_2675, f63);
and(x63, t_2674, t_2675);
not(t_2676, w59);
not(t_2677, g63);
and(y63, t_2676, t_2677);
not(t_2678, y61);
not(t_2679, g63);
and(z63, t_2678, t_2679);
not(t_2680, x62);
not(t_2681, h63);
and(a64, t_2680, t_2681);
not(t_2682, y62);
not(t_2683, i63);
and(b64, t_2682, t_2683);
not(t_2684, a63);
not(t_2685, j63);
and(c64, t_2684, t_2685);
not(t_2686, b63);
not(t_2687, s4);
and(d64, t_2686, t_2687);
not(t_2688, c63);
not(t_2689, k63);
and(e64, t_2688, t_2689);
not(t_2690, p62);
not(t_2691, i5);
and(f64, t_2690, t_2691);
not(t_2692, d63);
not(t_2693, l63);
and(g64, t_2692, t_2693);
not(t_2694, e63);
not(t_2695, m63);
and(h64, t_2694, t_2695);
not(t_2696, g63);
not(t_2697, v7);
and(i64, t_2696, t_2697);
not(t_2698, w62);
not(t_2699, l8);
and(j64, t_2698, t_2699);
not(t_2700, n63);
not(t_2701, o63);
and(k64, t_2700, t_2701);
not(t_2702, m62);
not(t_2703, p63);
and(l64, t_2702, t_2703);
not(t_2704, p63);
not(t_2705, n62);
and(m64, t_2704, t_2705);
not(t_2706, q63);
not(t_2707, r63);
and(n64, t_2706, t_2707);
not(t_2708, s63);
not(t_2709, d64);
and(o64, t_2708, t_2709);
not(t_2710, y60);
not(t_2711, f64);
and(p64, t_2710, t_2711);
not(t_2712, p62);
not(t_2713, f64);
and(q64, t_2712, t_2713);
not(t_2714, u63);
not(t_2715, v63);
and(r64, t_2714, t_2715);
not(t_2716, t62);
not(t_2717, w63);
and(s64, t_2716, t_2717);
not(t_2718, w63);
not(t_2719, u62);
and(t64, t_2718, t_2719);
not(t_2720, x63);
not(t_2721, y63);
and(u64, t_2720, t_2721);
not(t_2722, z63);
not(t_2723, i64);
and(v64, t_2722, t_2723);
not(t_2724, f61);
not(t_2725, j64);
and(w64, t_2724, t_2725);
not(t_2726, w62);
not(t_2727, j64);
and(x64, t_2726, t_2727);
not(t_2728, f64);
not(t_2729, i5);
and(y64, t_2728, t_2729);
not(t_2730, t63);
not(t_2731, y5);
and(z64, t_2730, t_2731);
not(t_2732, j64);
not(t_2733, l8);
and(a65, t_2732, t_2733);
not(t_2734, a64);
not(t_2735, b9);
and(b65, t_2734, t_2735);
not(t_2736, b64);
not(t_2737, r9);
and(c65, t_2736, t_2737);
not(t_2738, c64);
not(t_2739, h10);
and(d65, t_2738, t_2739);
not(t_2740, e64);
not(t_2741, x10);
and(e65, t_2740, t_2741);
not(t_2742, g64);
not(t_2743, n11);
and(f65, t_2742, t_2743);
not(t_2744, h64);
not(t_2745, d12);
and(g65, t_2744, t_2745);
not(t_2746, l64);
not(t_2747, m64);
and(h65, t_2746, t_2747);
not(t_2748, q63);
not(t_2749, n64);
and(i65, t_2748, t_2749);
not(t_2750, n64);
not(t_2751, r63);
and(j65, t_2750, t_2751);
not(t_2752, o64);
not(t_2753, p64);
and(k65, t_2752, t_2753);
not(t_2754, q64);
not(t_2755, y64);
and(l65, t_2754, t_2755);
not(t_2756, u61);
not(t_2757, z64);
and(m65, t_2756, t_2757);
not(t_2758, t63);
not(t_2759, z64);
and(n65, t_2758, t_2759);
not(t_2760, s64);
not(t_2761, t64);
and(o65, t_2760, t_2761);
not(t_2762, x63);
not(t_2763, u64);
and(p65, t_2762, t_2763);
not(t_2764, u64);
not(t_2765, y63);
and(q65, t_2764, t_2765);
not(t_2766, v64);
not(t_2767, w64);
and(r65, t_2766, t_2767);
not(t_2768, x64);
not(t_2769, a65);
and(s65, t_2768, t_2769);
not(t_2770, a64);
not(t_2771, b65);
and(t65, t_2770, t_2771);
not(t_2772, k64);
not(t_2773, l3);
and(u65, t_2772, t_2773);
not(t_2774, b64);
not(t_2775, c65);
and(v65, t_2774, t_2775);
not(t_2776, c64);
not(t_2777, d65);
and(w65, t_2776, t_2777);
not(t_2778, e64);
not(t_2779, e65);
and(x65, t_2778, t_2779);
not(t_2780, g64);
not(t_2781, f65);
and(y65, t_2780, t_2781);
not(t_2782, z64);
not(t_2783, y5);
and(z65, t_2782, t_2783);
not(t_2784, h64);
not(t_2785, g65);
and(a66, t_2784, t_2785);
not(t_2786, r64);
not(t_2787, o6);
and(b66, t_2786, t_2787);
not(t_2788, f62);
not(t_2789, b65);
and(c66, t_2788, t_2789);
not(t_2790, b65);
not(t_2791, b9);
and(d66, t_2790, t_2791);
not(t_2792, g62);
not(t_2793, c65);
and(e66, t_2792, t_2793);
not(t_2794, c65);
not(t_2795, r9);
and(f66, t_2794, t_2795);
not(t_2796, h62);
not(t_2797, d65);
and(g66, t_2796, t_2797);
not(t_2798, d65);
not(t_2799, h10);
and(h66, t_2798, t_2799);
not(t_2800, i62);
not(t_2801, e65);
and(i66, t_2800, t_2801);
not(t_2802, e65);
not(t_2803, x10);
and(j66, t_2802, t_2803);
not(t_2804, j62);
not(t_2805, f65);
and(k66, t_2804, t_2805);
not(t_2806, f65);
not(t_2807, n11);
and(l66, t_2806, t_2807);
not(t_2808, k62);
not(t_2809, g65);
and(m66, t_2808, t_2809);
not(t_2810, g65);
not(t_2811, d12);
and(n66, t_2810, t_2811);
not(t_2812, l62);
not(t_2813, u65);
and(o66, t_2812, t_2813);
not(t_2814, k64);
not(t_2815, u65);
and(p66, t_2814, t_2815);
not(t_2816, i65);
not(t_2817, j65);
and(q66, t_2816, t_2817);
not(t_2818, o64);
not(t_2819, k65);
and(r66, t_2818, t_2819);
not(t_2820, k65);
not(t_2821, p64);
and(s66, t_2820, t_2821);
not(t_2822, l65);
not(t_2823, m65);
and(t66, t_2822, t_2823);
not(t_2824, n65);
not(t_2825, z65);
and(u66, t_2824, t_2825);
not(t_2826, s62);
not(t_2827, b66);
and(v66, t_2826, t_2827);
not(t_2828, r64);
not(t_2829, b66);
and(w66, t_2828, t_2829);
not(t_2830, p65);
not(t_2831, q65);
and(x66, t_2830, t_2831);
not(t_2832, v64);
not(t_2833, r65);
and(y66, t_2832, t_2833);
not(t_2834, r65);
not(t_2835, w64);
and(z66, t_2834, t_2835);
not(t_2836, s65);
not(t_2837, c66);
and(a67, t_2836, t_2837);
not(t_2838, t65);
not(t_2839, d66);
and(b67, t_2838, t_2839);
not(t_2840, u65);
not(t_2841, l3);
and(c67, t_2840, t_2841);
not(t_2842, v65);
not(t_2843, f66);
and(d67, t_2842, t_2843);
not(t_2844, h65);
not(t_2845, b4);
and(e67, t_2844, t_2845);
not(t_2846, w65);
not(t_2847, h66);
and(f67, t_2846, t_2847);
not(t_2848, x65);
not(t_2849, j66);
and(g67, t_2848, t_2849);
not(t_2850, y65);
not(t_2851, l66);
and(h67, t_2850, t_2851);
not(t_2852, b66);
not(t_2853, o6);
and(i67, t_2852, t_2853);
not(t_2854, o65);
not(t_2855, e7);
and(j67, t_2854, t_2855);
not(t_2856, v2);
not(t_2857, o66);
and(k67, t_2856, t_2857);
not(t_2858, p66);
not(t_2859, c67);
and(l67, t_2858, t_2859);
not(t_2860, p63);
not(t_2861, e67);
and(m67, t_2860, t_2861);
not(t_2862, h65);
not(t_2863, e67);
and(n67, t_2862, t_2863);
not(t_2864, r66);
not(t_2865, s66);
and(o67, t_2864, t_2865);
not(t_2866, l65);
not(t_2867, t66);
and(p67, t_2866, t_2867);
not(t_2868, t66);
not(t_2869, m65);
and(q67, t_2868, t_2869);
not(t_2870, u66);
not(t_2871, v66);
and(r67, t_2870, t_2871);
not(t_2872, w66);
not(t_2873, i67);
and(s67, t_2872, t_2873);
not(t_2874, w63);
not(t_2875, j67);
and(t67, t_2874, t_2875);
not(t_2876, o65);
not(t_2877, j67);
and(u67, t_2876, t_2877);
not(t_2878, y66);
not(t_2879, z66);
and(v67, t_2878, t_2879);
not(t_2880, s65);
not(t_2881, a67);
and(w67, t_2880, t_2881);
not(t_2882, e67);
not(t_2883, b4);
and(x67, t_2882, t_2883);
not(t_2884, q66);
not(t_2885, r4);
and(y67, t_2884, t_2885);
not(t_2886, j67);
not(t_2887, e7);
and(z67, t_2886, t_2887);
not(t_2888, x66);
not(t_2889, u7);
and(a68, t_2888, t_2889);
not(t_2890, a67);
not(t_2891, c66);
and(b68, t_2890, t_2891);
not(t_2892, b67);
not(t_2893, e66);
and(c68, t_2892, t_2893);
not(t_2894, d67);
not(t_2895, g66);
and(d68, t_2894, t_2895);
not(t_2896, f67);
not(t_2897, i66);
and(e68, t_2896, t_2897);
not(t_2898, g67);
not(t_2899, k66);
and(f68, t_2898, t_2899);
not(t_2900, h67);
not(t_2901, m66);
and(g68, t_2900, t_2901);
not(t_2902, v2);
not(t_2903, k67);
and(h68, t_2902, t_2903);
not(t_2904, k67);
not(t_2905, o66);
and(i68, t_2904, t_2905);
not(t_2906, l67);
not(t_2907, m67);
and(j68, t_2906, t_2907);
not(t_2908, n67);
not(t_2909, x67);
and(k68, t_2908, t_2909);
not(t_2910, n64);
not(t_2911, y67);
and(l68, t_2910, t_2911);
not(t_2912, q66);
not(t_2913, y67);
and(m68, t_2912, t_2913);
not(t_2914, p67);
not(t_2915, q67);
and(n68, t_2914, t_2915);
not(t_2916, u66);
not(t_2917, r67);
and(o68, t_2916, t_2917);
not(t_2918, r67);
not(t_2919, v66);
and(p68, t_2918, t_2919);
not(t_2920, s67);
not(t_2921, t67);
and(q68, t_2920, t_2921);
not(t_2922, u67);
not(t_2923, z67);
and(r68, t_2922, t_2923);
not(t_2924, u64);
not(t_2925, a68);
and(s68, t_2924, t_2925);
not(t_2926, x66);
not(t_2927, a68);
and(t68, t_2926, t_2927);
not(t_2928, w67);
not(t_2929, b68);
and(u68, t_2928, t_2929);
not(t_2930, b67);
not(t_2931, c68);
and(v68, t_2930, t_2931);
not(t_2932, d67);
not(t_2933, d68);
and(w68, t_2932, t_2933);
not(t_2934, f67);
not(t_2935, e68);
and(x68, t_2934, t_2935);
not(t_2936, y67);
not(t_2937, r4);
and(y68, t_2936, t_2937);
not(t_2938, g67);
not(t_2939, f68);
and(z68, t_2938, t_2939);
not(t_2940, o67);
not(t_2941, h5);
and(a69, t_2940, t_2941);
not(t_2942, h67);
not(t_2943, g68);
and(b69, t_2942, t_2943);
not(t_2944, a68);
not(t_2945, u7);
and(c69, t_2944, t_2945);
not(t_2946, v67);
not(t_2947, k8);
and(d69, t_2946, t_2947);
not(t_2948, c68);
not(t_2949, e66);
and(e69, t_2948, t_2949);
not(t_2950, d68);
not(t_2951, g66);
and(f69, t_2950, t_2951);
not(t_2952, e68);
not(t_2953, i66);
and(g69, t_2952, t_2953);
not(t_2954, f68);
not(t_2955, k66);
and(h69, t_2954, t_2955);
not(t_2956, g68);
not(t_2957, m66);
and(i69, t_2956, t_2957);
not(t_2958, h68);
not(t_2959, i68);
and(j69, t_2958, t_2959);
not(t_2960, l67);
not(t_2961, j68);
and(k69, t_2960, t_2961);
not(t_2962, j68);
not(t_2963, m67);
and(l69, t_2962, t_2963);
not(t_2964, k68);
not(t_2965, l68);
and(m69, t_2964, t_2965);
not(t_2966, m68);
not(t_2967, y68);
and(n69, t_2966, t_2967);
not(t_2968, k65);
not(t_2969, a69);
and(o69, t_2968, t_2969);
not(t_2970, o67);
not(t_2971, a69);
and(p69, t_2970, t_2971);
not(t_2972, o68);
not(t_2973, p68);
and(q69, t_2972, t_2973);
not(t_2974, s67);
not(t_2975, q68);
and(r69, t_2974, t_2975);
not(t_2976, q68);
not(t_2977, t67);
and(s69, t_2976, t_2977);
not(t_2978, r68);
not(t_2979, s68);
and(t69, t_2978, t_2979);
not(t_2980, t68);
not(t_2981, c69);
and(u69, t_2980, t_2981);
not(t_2982, r65);
not(t_2983, d69);
and(v69, t_2982, t_2983);
not(t_2984, v67);
not(t_2985, d69);
and(w69, t_2984, t_2985);
not(t_2986, v68);
not(t_2987, e69);
and(x69, t_2986, t_2987);
not(t_2988, w68);
not(t_2989, f69);
and(y69, t_2988, t_2989);
not(t_2990, x68);
not(t_2991, g69);
and(z69, t_2990, t_2991);
not(t_2992, z68);
not(t_2993, h69);
and(a70, t_2992, t_2993);
not(t_2994, a69);
not(t_2995, h5);
and(b70, t_2994, t_2995);
not(t_2996, b69);
not(t_2997, i69);
and(c70, t_2996, t_2997);
not(t_2998, n68);
not(t_2999, x5);
and(d70, t_2998, t_2999);
not(t_3000, d69);
not(t_3001, k8);
and(e70, t_3000, t_3001);
not(t_3002, u68);
not(t_3003, a9);
and(f70, t_3002, t_3003);
not(t_3004, k69);
not(t_3005, l69);
and(g70, t_3004, t_3005);
not(t_3006, k68);
not(t_3007, m69);
and(h70, t_3006, t_3007);
not(t_3008, m69);
not(t_3009, l68);
and(i70, t_3008, t_3009);
not(t_3010, n69);
not(t_3011, o69);
and(j70, t_3010, t_3011);
not(t_3012, p69);
not(t_3013, b70);
and(k70, t_3012, t_3013);
not(t_3014, t66);
not(t_3015, d70);
and(l70, t_3014, t_3015);
not(t_3016, n68);
not(t_3017, d70);
and(m70, t_3016, t_3017);
not(t_3018, r69);
not(t_3019, s69);
and(n70, t_3018, t_3019);
not(t_3020, r68);
not(t_3021, t69);
and(o70, t_3020, t_3021);
not(t_3022, t69);
not(t_3023, s68);
and(p70, t_3022, t_3023);
not(t_3024, u69);
not(t_3025, v69);
and(q70, t_3024, t_3025);
not(t_3026, w69);
not(t_3027, e70);
and(r70, t_3026, t_3027);
not(t_3028, a67);
not(t_3029, f70);
and(s70, t_3028, t_3029);
not(t_3030, u68);
not(t_3031, f70);
and(t70, t_3030, t_3031);
not(t_3032, j69);
not(t_3033, k3);
and(u70, t_3032, t_3033);
not(t_3034, d70);
not(t_3035, x5);
and(v70, t_3034, t_3035);
not(t_3036, q69);
not(t_3037, n6);
and(w70, t_3036, t_3037);
not(t_3038, f70);
not(t_3039, a9);
and(x70, t_3038, t_3039);
not(t_3040, x69);
not(t_3041, q9);
and(y70, t_3040, t_3041);
not(t_3042, y69);
not(t_3043, g10);
and(z70, t_3042, t_3043);
not(t_3044, z69);
not(t_3045, w10);
and(a71, t_3044, t_3045);
not(t_3046, a70);
not(t_3047, m11);
and(b71, t_3046, t_3047);
not(t_3048, c70);
not(t_3049, c12);
and(c71, t_3048, t_3049);
not(t_3050, k67);
not(t_3051, u70);
and(d71, t_3050, t_3051);
not(t_3052, j69);
not(t_3053, u70);
and(e71, t_3052, t_3053);
not(t_3054, h70);
not(t_3055, i70);
and(f71, t_3054, t_3055);
not(t_3056, n69);
not(t_3057, j70);
and(g71, t_3056, t_3057);
not(t_3058, j70);
not(t_3059, o69);
and(h71, t_3058, t_3059);
not(t_3060, k70);
not(t_3061, l70);
and(i71, t_3060, t_3061);
not(t_3062, m70);
not(t_3063, v70);
and(j71, t_3062, t_3063);
not(t_3064, r67);
not(t_3065, w70);
and(k71, t_3064, t_3065);
not(t_3066, q69);
not(t_3067, w70);
and(l71, t_3066, t_3067);
not(t_3068, o70);
not(t_3069, p70);
and(m71, t_3068, t_3069);
not(t_3070, u69);
not(t_3071, q70);
and(n71, t_3070, t_3071);
not(t_3072, q70);
not(t_3073, v69);
and(o71, t_3072, t_3073);
not(t_3074, r70);
not(t_3075, s70);
and(p71, t_3074, t_3075);
not(t_3076, t70);
not(t_3077, x70);
and(q71, t_3076, t_3077);
not(t_3078, x69);
not(t_3079, y70);
and(r71, t_3078, t_3079);
not(t_3080, u70);
not(t_3081, k3);
and(s71, t_3080, t_3081);
not(t_3082, y69);
not(t_3083, z70);
and(t71, t_3082, t_3083);
not(t_3084, g70);
not(t_3085, a4);
and(u71, t_3084, t_3085);
not(t_3086, z69);
not(t_3087, a71);
and(v71, t_3086, t_3087);
not(t_3088, a70);
not(t_3089, b71);
and(w71, t_3088, t_3089);
not(t_3090, c70);
not(t_3091, c71);
and(x71, t_3090, t_3091);
not(t_3092, w70);
not(t_3093, n6);
and(y71, t_3092, t_3093);
not(t_3094, n70);
not(t_3095, d7);
and(z71, t_3094, t_3095);
not(t_3096, c68);
not(t_3097, y70);
and(a72, t_3096, t_3097);
not(t_3098, y70);
not(t_3099, q9);
and(b72, t_3098, t_3099);
not(t_3100, d68);
not(t_3101, z70);
and(c72, t_3100, t_3101);
not(t_3102, z70);
not(t_3103, g10);
and(d72, t_3102, t_3103);
not(t_3104, e68);
not(t_3105, a71);
and(e72, t_3104, t_3105);
not(t_3106, a71);
not(t_3107, w10);
and(f72, t_3106, t_3107);
not(t_3108, f68);
not(t_3109, b71);
and(g72, t_3108, t_3109);
not(t_3110, b71);
not(t_3111, m11);
and(h72, t_3110, t_3111);
not(t_3112, g68);
not(t_3113, c71);
and(i72, t_3112, t_3113);
not(t_3114, c71);
not(t_3115, c12);
and(j72, t_3114, t_3115);
not(t_3116, u2);
not(t_3117, d71);
and(k72, t_3116, t_3117);
not(t_3118, e71);
not(t_3119, s71);
and(l72, t_3118, t_3119);
not(t_3120, j68);
not(t_3121, u71);
and(m72, t_3120, t_3121);
not(t_3122, g70);
not(t_3123, u71);
and(n72, t_3122, t_3123);
not(t_3124, g71);
not(t_3125, h71);
and(o72, t_3124, t_3125);
not(t_3126, k70);
not(t_3127, i71);
and(p72, t_3126, t_3127);
not(t_3128, i71);
not(t_3129, l70);
and(q72, t_3128, t_3129);
not(t_3130, j71);
not(t_3131, k71);
and(r72, t_3130, t_3131);
not(t_3132, l71);
not(t_3133, y71);
and(s72, t_3132, t_3133);
not(t_3134, q68);
not(t_3135, z71);
and(t72, t_3134, t_3135);
not(t_3136, n70);
not(t_3137, z71);
and(u72, t_3136, t_3137);
not(t_3138, n71);
not(t_3139, o71);
and(v72, t_3138, t_3139);
not(t_3140, r70);
not(t_3141, p71);
and(w72, t_3140, t_3141);
not(t_3142, p71);
not(t_3143, s70);
and(x72, t_3142, t_3143);
not(t_3144, q71);
not(t_3145, a72);
and(y72, t_3144, t_3145);
not(t_3146, r71);
not(t_3147, b72);
and(z72, t_3146, t_3147);
not(t_3148, t71);
not(t_3149, d72);
and(a73, t_3148, t_3149);
not(t_3150, u71);
not(t_3151, a4);
and(b73, t_3150, t_3151);
not(t_3152, v71);
not(t_3153, f72);
and(c73, t_3152, t_3153);
not(t_3154, f71);
not(t_3155, q4);
and(d73, t_3154, t_3155);
not(t_3156, w71);
not(t_3157, h72);
and(e73, t_3156, t_3157);
not(t_3158, z71);
not(t_3159, d7);
and(f73, t_3158, t_3159);
not(t_3160, m71);
not(t_3161, t7);
and(g73, t_3160, t_3161);
not(t_3162, u2);
not(t_3163, k72);
and(h73, t_3162, t_3163);
not(t_3164, k72);
not(t_3165, d71);
and(i73, t_3164, t_3165);
not(t_3166, l72);
not(t_3167, m72);
and(j73, t_3166, t_3167);
not(t_3168, n72);
not(t_3169, b73);
and(k73, t_3168, t_3169);
not(t_3170, m69);
not(t_3171, d73);
and(l73, t_3170, t_3171);
not(t_3172, f71);
not(t_3173, d73);
and(m73, t_3172, t_3173);
not(t_3174, p72);
not(t_3175, q72);
and(n73, t_3174, t_3175);
not(t_3176, j71);
not(t_3177, r72);
and(o73, t_3176, t_3177);
not(t_3178, r72);
not(t_3179, k71);
and(p73, t_3178, t_3179);
not(t_3180, s72);
not(t_3181, t72);
and(q73, t_3180, t_3181);
not(t_3182, u72);
not(t_3183, f73);
and(r73, t_3182, t_3183);
not(t_3184, t69);
not(t_3185, g73);
and(s73, t_3184, t_3185);
not(t_3186, m71);
not(t_3187, g73);
and(t73, t_3186, t_3187);
not(t_3188, w72);
not(t_3189, x72);
and(u73, t_3188, t_3189);
not(t_3190, q71);
not(t_3191, y72);
and(v73, t_3190, t_3191);
not(t_3192, d73);
not(t_3193, q4);
and(w73, t_3192, t_3193);
not(t_3194, o72);
not(t_3195, g5);
and(x73, t_3194, t_3195);
not(t_3196, g73);
not(t_3197, t7);
and(y73, t_3196, t_3197);
not(t_3198, v72);
not(t_3199, j8);
and(z73, t_3198, t_3199);
not(t_3200, y72);
not(t_3201, a72);
and(a74, t_3200, t_3201);
not(t_3202, z72);
not(t_3203, c72);
and(b74, t_3202, t_3203);
not(t_3204, a73);
not(t_3205, e72);
and(c74, t_3204, t_3205);
not(t_3206, c73);
not(t_3207, g72);
and(d74, t_3206, t_3207);
not(t_3208, e73);
not(t_3209, i72);
and(e74, t_3208, t_3209);
not(t_3210, h73);
not(t_3211, i73);
and(f74, t_3210, t_3211);
not(t_3212, l72);
not(t_3213, j73);
and(g74, t_3212, t_3213);
not(t_3214, j73);
not(t_3215, m72);
and(h74, t_3214, t_3215);
not(t_3216, k73);
not(t_3217, l73);
and(i74, t_3216, t_3217);
not(t_3218, m73);
not(t_3219, w73);
and(j74, t_3218, t_3219);
not(t_3220, j70);
not(t_3221, x73);
and(k74, t_3220, t_3221);
not(t_3222, o72);
not(t_3223, x73);
and(l74, t_3222, t_3223);
not(t_3224, o73);
not(t_3225, p73);
and(m74, t_3224, t_3225);
not(t_3226, s72);
not(t_3227, q73);
and(n74, t_3226, t_3227);
not(t_3228, q73);
not(t_3229, t72);
and(o74, t_3228, t_3229);
not(t_3230, r73);
not(t_3231, s73);
and(p74, t_3230, t_3231);
not(t_3232, t73);
not(t_3233, y73);
and(q74, t_3232, t_3233);
not(t_3234, q70);
not(t_3235, z73);
and(r74, t_3234, t_3235);
not(t_3236, v72);
not(t_3237, z73);
and(s74, t_3236, t_3237);
not(t_3238, v73);
not(t_3239, a74);
and(t74, t_3238, t_3239);
not(t_3240, z72);
not(t_3241, b74);
and(u74, t_3240, t_3241);
not(t_3242, a73);
not(t_3243, c74);
and(v74, t_3242, t_3243);
not(t_3244, c73);
not(t_3245, d74);
and(w74, t_3244, t_3245);
not(t_3246, e73);
not(t_3247, e74);
and(x74, t_3246, t_3247);
not(t_3248, x73);
not(t_3249, g5);
and(y74, t_3248, t_3249);
not(t_3250, n73);
not(t_3251, w5);
and(z74, t_3250, t_3251);
not(t_3252, z73);
not(t_3253, j8);
and(a75, t_3252, t_3253);
not(t_3254, u73);
not(t_3255, z8);
and(b75, t_3254, t_3255);
not(t_3256, b74);
not(t_3257, c72);
and(c75, t_3256, t_3257);
not(t_3258, c74);
not(t_3259, e72);
and(d75, t_3258, t_3259);
not(t_3260, d74);
not(t_3261, g72);
and(e75, t_3260, t_3261);
not(t_3262, e74);
not(t_3263, i72);
and(f75, t_3262, t_3263);
not(t_3264, g74);
not(t_3265, h74);
and(g75, t_3264, t_3265);
not(t_3266, k73);
not(t_3267, i74);
and(h75, t_3266, t_3267);
not(t_3268, i74);
not(t_3269, l73);
and(i75, t_3268, t_3269);
not(t_3270, j74);
not(t_3271, k74);
and(j75, t_3270, t_3271);
not(t_3272, l74);
not(t_3273, y74);
and(k75, t_3272, t_3273);
not(t_3274, i71);
not(t_3275, z74);
and(l75, t_3274, t_3275);
not(t_3276, n73);
not(t_3277, z74);
and(m75, t_3276, t_3277);
not(t_3278, n74);
not(t_3279, o74);
and(n75, t_3278, t_3279);
not(t_3280, r73);
not(t_3281, p74);
and(o75, t_3280, t_3281);
not(t_3282, p74);
not(t_3283, s73);
and(p75, t_3282, t_3283);
not(t_3284, q74);
not(t_3285, r74);
and(q75, t_3284, t_3285);
not(t_3286, s74);
not(t_3287, a75);
and(r75, t_3286, t_3287);
not(t_3288, p71);
not(t_3289, b75);
and(s75, t_3288, t_3289);
not(t_3290, u73);
not(t_3291, b75);
and(t75, t_3290, t_3291);
not(t_3292, u74);
not(t_3293, c75);
and(u75, t_3292, t_3293);
not(t_3294, f74);
not(t_3295, j3);
and(v75, t_3294, t_3295);
not(t_3296, v74);
not(t_3297, d75);
and(w75, t_3296, t_3297);
not(t_3298, w74);
not(t_3299, e75);
and(x75, t_3298, t_3299);
not(t_3300, x74);
not(t_3301, f75);
and(y75, t_3300, t_3301);
not(t_3302, z74);
not(t_3303, w5);
and(z75, t_3302, t_3303);
not(t_3304, m74);
not(t_3305, m6);
and(a76, t_3304, t_3305);
not(t_3306, b75);
not(t_3307, z8);
and(b76, t_3306, t_3307);
not(t_3308, t74);
not(t_3309, p9);
and(c76, t_3308, t_3309);
not(t_3310, k72);
not(t_3311, v75);
and(d76, t_3310, t_3311);
not(t_3312, f74);
not(t_3313, v75);
and(e76, t_3312, t_3313);
not(t_3314, h75);
not(t_3315, i75);
and(f76, t_3314, t_3315);
not(t_3316, j74);
not(t_3317, j75);
and(g76, t_3316, t_3317);
not(t_3318, j75);
not(t_3319, k74);
and(h76, t_3318, t_3319);
not(t_3320, k75);
not(t_3321, l75);
and(i76, t_3320, t_3321);
not(t_3322, m75);
not(t_3323, z75);
and(j76, t_3322, t_3323);
not(t_3324, r72);
not(t_3325, a76);
and(k76, t_3324, t_3325);
not(t_3326, m74);
not(t_3327, a76);
and(l76, t_3326, t_3327);
not(t_3328, o75);
not(t_3329, p75);
and(m76, t_3328, t_3329);
not(t_3330, q74);
not(t_3331, q75);
and(n76, t_3330, t_3331);
not(t_3332, q75);
not(t_3333, r74);
and(o76, t_3332, t_3333);
not(t_3334, r75);
not(t_3335, s75);
and(p76, t_3334, t_3335);
not(t_3336, t75);
not(t_3337, b76);
and(q76, t_3336, t_3337);
not(t_3338, y72);
not(t_3339, c76);
and(r76, t_3338, t_3339);
not(t_3340, t74);
not(t_3341, c76);
and(s76, t_3340, t_3341);
not(t_3342, v75);
not(t_3343, j3);
and(t76, t_3342, t_3343);
not(t_3344, g75);
not(t_3345, z3);
and(u76, t_3344, t_3345);
not(t_3346, a76);
not(t_3347, m6);
and(v76, t_3346, t_3347);
not(t_3348, n75);
not(t_3349, c7);
and(w76, t_3348, t_3349);
not(t_3350, c76);
not(t_3351, p9);
and(x76, t_3350, t_3351);
not(t_3352, u75);
not(t_3353, f10);
and(y76, t_3352, t_3353);
not(t_3354, w75);
not(t_3355, v10);
and(z76, t_3354, t_3355);
not(t_3356, x75);
not(t_3357, l11);
and(a77, t_3356, t_3357);
not(t_3358, y75);
not(t_3359, b12);
and(b77, t_3358, t_3359);
not(t_3360, t2);
not(t_3361, d76);
and(c77, t_3360, t_3361);
not(t_3362, e76);
not(t_3363, t76);
and(d77, t_3362, t_3363);
not(t_3364, j73);
not(t_3365, u76);
and(e77, t_3364, t_3365);
not(t_3366, g75);
not(t_3367, u76);
and(f77, t_3366, t_3367);
not(t_3368, g76);
not(t_3369, h76);
and(g77, t_3368, t_3369);
not(t_3370, k75);
not(t_3371, i76);
and(h77, t_3370, t_3371);
not(t_3372, i76);
not(t_3373, l75);
and(i77, t_3372, t_3373);
not(t_3374, j76);
not(t_3375, k76);
and(j77, t_3374, t_3375);
not(t_3376, l76);
not(t_3377, v76);
and(k77, t_3376, t_3377);
not(t_3378, q73);
not(t_3379, w76);
and(l77, t_3378, t_3379);
not(t_3380, n75);
not(t_3381, w76);
and(m77, t_3380, t_3381);
not(t_3382, n76);
not(t_3383, o76);
and(n77, t_3382, t_3383);
not(t_3384, r75);
not(t_3385, p76);
and(o77, t_3384, t_3385);
not(t_3386, p76);
not(t_3387, s75);
and(p77, t_3386, t_3387);
not(t_3388, q76);
not(t_3389, r76);
and(q77, t_3388, t_3389);
not(t_3390, s76);
not(t_3391, x76);
and(r77, t_3390, t_3391);
not(t_3392, u75);
not(t_3393, y76);
and(s77, t_3392, t_3393);
not(t_3394, w75);
not(t_3395, z76);
and(t77, t_3394, t_3395);
not(t_3396, u76);
not(t_3397, z3);
and(u77, t_3396, t_3397);
not(t_3398, x75);
not(t_3399, a77);
and(v77, t_3398, t_3399);
not(t_3400, f76);
not(t_3401, p4);
and(w77, t_3400, t_3401);
not(t_3402, y75);
not(t_3403, b77);
and(x77, t_3402, t_3403);
not(t_3404, w76);
not(t_3405, c7);
and(y77, t_3404, t_3405);
not(t_3406, m76);
not(t_3407, s7);
and(z77, t_3406, t_3407);
not(t_3408, b74);
not(t_3409, y76);
and(a78, t_3408, t_3409);
not(t_3410, y76);
not(t_3411, f10);
and(b78, t_3410, t_3411);
not(t_3412, c74);
not(t_3413, z76);
and(c78, t_3412, t_3413);
not(t_3414, z76);
not(t_3415, v10);
and(d78, t_3414, t_3415);
not(t_3416, d74);
not(t_3417, a77);
and(e78, t_3416, t_3417);
not(t_3418, a77);
not(t_3419, l11);
and(f78, t_3418, t_3419);
not(t_3420, e74);
not(t_3421, b77);
and(g78, t_3420, t_3421);
not(t_3422, b77);
not(t_3423, b12);
and(h78, t_3422, t_3423);
not(t_3424, t2);
not(t_3425, c77);
and(i78, t_3424, t_3425);
not(t_3426, c77);
not(t_3427, d76);
and(j78, t_3426, t_3427);
not(t_3428, d77);
not(t_3429, e77);
and(k78, t_3428, t_3429);
not(t_3430, f77);
not(t_3431, u77);
and(l78, t_3430, t_3431);
not(t_3432, i74);
not(t_3433, w77);
and(m78, t_3432, t_3433);
not(t_3434, f76);
not(t_3435, w77);
and(n78, t_3434, t_3435);
not(t_3436, h77);
not(t_3437, i77);
and(o78, t_3436, t_3437);
not(t_3438, j76);
not(t_3439, j77);
and(p78, t_3438, t_3439);
not(t_3440, j77);
not(t_3441, k76);
and(q78, t_3440, t_3441);
not(t_3442, k77);
not(t_3443, l77);
and(r78, t_3442, t_3443);
not(t_3444, m77);
not(t_3445, y77);
and(s78, t_3444, t_3445);
not(t_3446, p74);
not(t_3447, z77);
and(t78, t_3446, t_3447);
not(t_3448, m76);
not(t_3449, z77);
and(u78, t_3448, t_3449);
not(t_3450, o77);
not(t_3451, p77);
and(v78, t_3450, t_3451);
not(t_3452, q76);
not(t_3453, q77);
and(w78, t_3452, t_3453);
not(t_3454, q77);
not(t_3455, r76);
and(x78, t_3454, t_3455);
not(t_3456, r77);
not(t_3457, a78);
and(y78, t_3456, t_3457);
not(t_3458, s77);
not(t_3459, b78);
and(z78, t_3458, t_3459);
not(t_3460, t77);
not(t_3461, d78);
and(a79, t_3460, t_3461);
not(t_3462, v77);
not(t_3463, f78);
and(b79, t_3462, t_3463);
not(t_3464, w77);
not(t_3465, p4);
and(c79, t_3464, t_3465);
not(t_3466, g77);
not(t_3467, f5);
and(d79, t_3466, t_3467);
not(t_3468, z77);
not(t_3469, s7);
and(e79, t_3468, t_3469);
not(t_3470, n77);
not(t_3471, i8);
and(f79, t_3470, t_3471);
not(t_3472, i78);
not(t_3473, j78);
and(g79, t_3472, t_3473);
not(t_3474, d77);
not(t_3475, k78);
and(h79, t_3474, t_3475);
not(t_3476, k78);
not(t_3477, e77);
and(i79, t_3476, t_3477);
not(t_3478, l78);
not(t_3479, m78);
and(j79, t_3478, t_3479);
not(t_3480, n78);
not(t_3481, c79);
and(k79, t_3480, t_3481);
not(t_3482, j75);
not(t_3483, d79);
and(l79, t_3482, t_3483);
not(t_3484, g77);
not(t_3485, d79);
and(m79, t_3484, t_3485);
not(t_3486, p78);
not(t_3487, q78);
and(n79, t_3486, t_3487);
not(t_3488, k77);
not(t_3489, r78);
and(o79, t_3488, t_3489);
not(t_3490, r78);
not(t_3491, l77);
and(p79, t_3490, t_3491);
not(t_3492, s78);
not(t_3493, t78);
and(q79, t_3492, t_3493);
not(t_3494, u78);
not(t_3495, e79);
and(r79, t_3494, t_3495);
not(t_3496, q75);
not(t_3497, f79);
and(s79, t_3496, t_3497);
not(t_3498, n77);
not(t_3499, f79);
and(t79, t_3498, t_3499);
not(t_3500, w78);
not(t_3501, x78);
and(u79, t_3500, t_3501);
not(t_3502, r77);
not(t_3503, y78);
and(v79, t_3502, t_3503);
not(t_3504, d79);
not(t_3505, f5);
and(w79, t_3504, t_3505);
not(t_3506, o78);
not(t_3507, v5);
and(x79, t_3506, t_3507);
not(t_3508, f79);
not(t_3509, i8);
and(y79, t_3508, t_3509);
not(t_3510, v78);
not(t_3511, y8);
and(z79, t_3510, t_3511);
not(t_3512, y78);
not(t_3513, a78);
and(a80, t_3512, t_3513);
not(t_3514, z78);
not(t_3515, c78);
and(b80, t_3514, t_3515);
not(t_3516, a79);
not(t_3517, e78);
and(c80, t_3516, t_3517);
not(t_3518, b79);
not(t_3519, g78);
and(d80, t_3518, t_3519);
not(t_3520, h79);
not(t_3521, i79);
and(e80, t_3520, t_3521);
not(t_3522, l78);
not(t_3523, j79);
and(f80, t_3522, t_3523);
not(t_3524, j79);
not(t_3525, m78);
and(g80, t_3524, t_3525);
not(t_3526, k79);
not(t_3527, l79);
and(h80, t_3526, t_3527);
not(t_3528, m79);
not(t_3529, w79);
and(i80, t_3528, t_3529);
not(t_3530, i76);
not(t_3531, x79);
and(j80, t_3530, t_3531);
not(t_3532, o78);
not(t_3533, x79);
and(k80, t_3532, t_3533);
not(t_3534, o79);
not(t_3535, p79);
and(l80, t_3534, t_3535);
not(t_3536, s78);
not(t_3537, q79);
and(m80, t_3536, t_3537);
not(t_3538, q79);
not(t_3539, t78);
and(n80, t_3538, t_3539);
not(t_3540, r79);
not(t_3541, s79);
and(o80, t_3540, t_3541);
not(t_3542, t79);
not(t_3543, y79);
and(p80, t_3542, t_3543);
not(t_3544, p76);
not(t_3545, z79);
and(q80, t_3544, t_3545);
not(t_3546, v78);
not(t_3547, z79);
and(r80, t_3546, t_3547);
not(t_3548, v79);
not(t_3549, a80);
and(s80, t_3548, t_3549);
not(t_3550, z78);
not(t_3551, b80);
and(t80, t_3550, t_3551);
not(t_3552, g79);
not(t_3553, i3);
and(u80, t_3552, t_3553);
not(t_3554, a79);
not(t_3555, c80);
and(v80, t_3554, t_3555);
not(t_3556, b79);
not(t_3557, d80);
and(w80, t_3556, t_3557);
not(t_3558, x79);
not(t_3559, v5);
and(x80, t_3558, t_3559);
not(t_3560, n79);
not(t_3561, l6);
and(y80, t_3560, t_3561);
not(t_3562, z79);
not(t_3563, y8);
and(z80, t_3562, t_3563);
not(t_3564, u79);
not(t_3565, o9);
and(a81, t_3564, t_3565);
not(t_3566, b80);
not(t_3567, c78);
and(b81, t_3566, t_3567);
not(t_3568, c80);
not(t_3569, e78);
and(c81, t_3568, t_3569);
not(t_3570, d80);
not(t_3571, g78);
and(d81, t_3570, t_3571);
not(t_3572, c77);
not(t_3573, u80);
and(e81, t_3572, t_3573);
not(t_3574, g79);
not(t_3575, u80);
and(f81, t_3574, t_3575);
not(t_3576, f80);
not(t_3577, g80);
and(g81, t_3576, t_3577);
not(t_3578, k79);
not(t_3579, h80);
and(h81, t_3578, t_3579);
not(t_3580, h80);
not(t_3581, l79);
and(i81, t_3580, t_3581);
not(t_3582, i80);
not(t_3583, j80);
and(j81, t_3582, t_3583);
not(t_3584, k80);
not(t_3585, x80);
and(k81, t_3584, t_3585);
not(t_3586, j77);
not(t_3587, y80);
and(l81, t_3586, t_3587);
not(t_3588, n79);
not(t_3589, y80);
and(m81, t_3588, t_3589);
not(t_3590, m80);
not(t_3591, n80);
and(n81, t_3590, t_3591);
not(t_3592, r79);
not(t_3593, o80);
and(o81, t_3592, t_3593);
not(t_3594, o80);
not(t_3595, s79);
and(p81, t_3594, t_3595);
not(t_3596, p80);
not(t_3597, q80);
and(q81, t_3596, t_3597);
not(t_3598, r80);
not(t_3599, z80);
and(r81, t_3598, t_3599);
not(t_3600, q77);
not(t_3601, a81);
and(s81, t_3600, t_3601);
not(t_3602, u79);
not(t_3603, a81);
and(t81, t_3602, t_3603);
not(t_3604, t80);
not(t_3605, b81);
and(u81, t_3604, t_3605);
not(t_3606, u80);
not(t_3607, i3);
and(v81, t_3606, t_3607);
not(t_3608, v80);
not(t_3609, c81);
and(w81, t_3608, t_3609);
not(t_3610, e80);
not(t_3611, y3);
and(x81, t_3610, t_3611);
not(t_3612, w80);
not(t_3613, d81);
and(y81, t_3612, t_3613);
not(t_3614, y80);
not(t_3615, l6);
and(z81, t_3614, t_3615);
not(t_3616, l80);
not(t_3617, b7);
and(a82, t_3616, t_3617);
not(t_3618, a81);
not(t_3619, o9);
and(b82, t_3618, t_3619);
not(t_3620, s80);
not(t_3621, e10);
and(c82, t_3620, t_3621);
not(t_3622, s2);
not(t_3623, e81);
and(d82, t_3622, t_3623);
not(t_3624, f81);
not(t_3625, v81);
and(e82, t_3624, t_3625);
not(t_3626, k78);
not(t_3627, x81);
and(f82, t_3626, t_3627);
not(t_3628, e80);
not(t_3629, x81);
and(g82, t_3628, t_3629);
not(t_3630, h81);
not(t_3631, i81);
and(h82, t_3630, t_3631);
not(t_3632, i80);
not(t_3633, j81);
and(i82, t_3632, t_3633);
not(t_3634, j81);
not(t_3635, j80);
and(j82, t_3634, t_3635);
not(t_3636, k81);
not(t_3637, l81);
and(k82, t_3636, t_3637);
not(t_3638, m81);
not(t_3639, z81);
and(l82, t_3638, t_3639);
not(t_3640, r78);
not(t_3641, a82);
and(m82, t_3640, t_3641);
not(t_3642, l80);
not(t_3643, a82);
and(n82, t_3642, t_3643);
not(t_3644, o81);
not(t_3645, p81);
and(o82, t_3644, t_3645);
not(t_3646, p80);
not(t_3647, q81);
and(p82, t_3646, t_3647);
not(t_3648, q81);
not(t_3649, q80);
and(q82, t_3648, t_3649);
not(t_3650, r81);
not(t_3651, s81);
and(r82, t_3650, t_3651);
not(t_3652, t81);
not(t_3653, b82);
and(s82, t_3652, t_3653);
not(t_3654, y78);
not(t_3655, c82);
and(t82, t_3654, t_3655);
not(t_3656, s80);
not(t_3657, c82);
and(u82, t_3656, t_3657);
not(t_3658, x81);
not(t_3659, y3);
and(v82, t_3658, t_3659);
not(t_3660, g81);
not(t_3661, o4);
and(w82, t_3660, t_3661);
not(t_3662, a82);
not(t_3663, b7);
and(x82, t_3662, t_3663);
not(t_3664, n81);
not(t_3665, r7);
and(y82, t_3664, t_3665);
not(t_3666, c82);
not(t_3667, e10);
and(z82, t_3666, t_3667);
not(t_3668, u81);
not(t_3669, u10);
and(a83, t_3668, t_3669);
not(t_3670, w81);
not(t_3671, k11);
and(b83, t_3670, t_3671);
not(t_3672, y81);
not(t_3673, a12);
and(c83, t_3672, t_3673);
not(t_3674, s2);
not(t_3675, d82);
and(d83, t_3674, t_3675);
not(t_3676, d82);
not(t_3677, e81);
and(e83, t_3676, t_3677);
not(t_3678, e82);
not(t_3679, f82);
and(f83, t_3678, t_3679);
not(t_3680, g82);
not(t_3681, v82);
and(g83, t_3680, t_3681);
not(t_3682, j79);
not(t_3683, w82);
and(h83, t_3682, t_3683);
not(t_3684, g81);
not(t_3685, w82);
and(i83, t_3684, t_3685);
not(t_3686, i82);
not(t_3687, j82);
and(j83, t_3686, t_3687);
not(t_3688, k81);
not(t_3689, k82);
and(k83, t_3688, t_3689);
not(t_3690, k82);
not(t_3691, l81);
and(l83, t_3690, t_3691);
not(t_3692, l82);
not(t_3693, m82);
and(m83, t_3692, t_3693);
not(t_3694, n82);
not(t_3695, x82);
and(n83, t_3694, t_3695);
not(t_3696, q79);
not(t_3697, y82);
and(o83, t_3696, t_3697);
not(t_3698, n81);
not(t_3699, y82);
and(p83, t_3698, t_3699);
not(t_3700, p82);
not(t_3701, q82);
and(q83, t_3700, t_3701);
not(t_3702, r81);
not(t_3703, r82);
and(r83, t_3702, t_3703);
not(t_3704, r82);
not(t_3705, s81);
and(s83, t_3704, t_3705);
not(t_3706, s82);
not(t_3707, t82);
and(t83, t_3706, t_3707);
not(t_3708, u82);
not(t_3709, z82);
and(u83, t_3708, t_3709);
not(t_3710, u81);
not(t_3711, a83);
and(v83, t_3710, t_3711);
not(t_3712, w81);
not(t_3713, b83);
and(w83, t_3712, t_3713);
not(t_3714, y81);
not(t_3715, c83);
and(x83, t_3714, t_3715);
not(t_3716, w82);
not(t_3717, o4);
and(y83, t_3716, t_3717);
not(t_3718, h82);
not(t_3719, e5);
and(z83, t_3718, t_3719);
not(t_3720, y82);
not(t_3721, r7);
and(a84, t_3720, t_3721);
not(t_3722, o82);
not(t_3723, h8);
and(b84, t_3722, t_3723);
not(t_3724, b80);
not(t_3725, a83);
and(c84, t_3724, t_3725);
not(t_3726, a83);
not(t_3727, u10);
and(d84, t_3726, t_3727);
not(t_3728, c80);
not(t_3729, b83);
and(e84, t_3728, t_3729);
not(t_3730, b83);
not(t_3731, k11);
and(f84, t_3730, t_3731);
not(t_3732, d80);
not(t_3733, c83);
and(g84, t_3732, t_3733);
not(t_3734, c83);
not(t_3735, a12);
and(h84, t_3734, t_3735);
not(t_3736, d83);
not(t_3737, e83);
and(i84, t_3736, t_3737);
not(t_3738, e82);
not(t_3739, f83);
and(j84, t_3738, t_3739);
not(t_3740, f83);
not(t_3741, f82);
and(k84, t_3740, t_3741);
not(t_3742, g83);
not(t_3743, h83);
and(l84, t_3742, t_3743);
not(t_3744, i83);
not(t_3745, y83);
and(m84, t_3744, t_3745);
not(t_3746, h80);
not(t_3747, z83);
and(n84, t_3746, t_3747);
not(t_3748, h82);
not(t_3749, z83);
and(o84, t_3748, t_3749);
not(t_3750, k83);
not(t_3751, l83);
and(p84, t_3750, t_3751);
not(t_3752, l82);
not(t_3753, m83);
and(q84, t_3752, t_3753);
not(t_3754, m83);
not(t_3755, m82);
and(r84, t_3754, t_3755);
not(t_3756, n83);
not(t_3757, o83);
and(s84, t_3756, t_3757);
not(t_3758, p83);
not(t_3759, a84);
and(t84, t_3758, t_3759);
not(t_3760, o80);
not(t_3761, b84);
and(u84, t_3760, t_3761);
not(t_3762, o82);
not(t_3763, b84);
and(v84, t_3762, t_3763);
not(t_3764, r83);
not(t_3765, s83);
and(w84, t_3764, t_3765);
not(t_3766, s82);
not(t_3767, t83);
and(x84, t_3766, t_3767);
not(t_3768, t83);
not(t_3769, t82);
and(y84, t_3768, t_3769);
not(t_3770, u83);
not(t_3771, c84);
and(z84, t_3770, t_3771);
not(t_3772, v83);
not(t_3773, d84);
and(a85, t_3772, t_3773);
not(t_3774, w83);
not(t_3775, f84);
and(b85, t_3774, t_3775);
not(t_3776, z83);
not(t_3777, e5);
and(c85, t_3776, t_3777);
not(t_3778, j83);
not(t_3779, u5);
and(d85, t_3778, t_3779);
not(t_3780, b84);
not(t_3781, h8);
and(e85, t_3780, t_3781);
not(t_3782, q83);
not(t_3783, x8);
and(f85, t_3782, t_3783);
not(t_3784, j84);
not(t_3785, k84);
and(g85, t_3784, t_3785);
not(t_3786, g83);
not(t_3787, l84);
and(h85, t_3786, t_3787);
not(t_3788, l84);
not(t_3789, h83);
and(i85, t_3788, t_3789);
not(t_3790, m84);
not(t_3791, n84);
and(j85, t_3790, t_3791);
not(t_3792, o84);
not(t_3793, c85);
and(k85, t_3792, t_3793);
not(t_3794, j81);
not(t_3795, d85);
and(l85, t_3794, t_3795);
not(t_3796, j83);
not(t_3797, d85);
and(m85, t_3796, t_3797);
not(t_3798, q84);
not(t_3799, r84);
and(n85, t_3798, t_3799);
not(t_3800, n83);
not(t_3801, s84);
and(o85, t_3800, t_3801);
not(t_3802, s84);
not(t_3803, o83);
and(p85, t_3802, t_3803);
not(t_3804, t84);
not(t_3805, u84);
and(q85, t_3804, t_3805);
not(t_3806, v84);
not(t_3807, e85);
and(r85, t_3806, t_3807);
not(t_3808, q81);
not(t_3809, f85);
and(s85, t_3808, t_3809);
not(t_3810, q83);
not(t_3811, f85);
and(t85, t_3810, t_3811);
not(t_3812, x84);
not(t_3813, y84);
and(u85, t_3812, t_3813);
not(t_3814, u83);
not(t_3815, z84);
and(v85, t_3814, t_3815);
not(t_3816, d85);
not(t_3817, u5);
and(w85, t_3816, t_3817);
not(t_3818, p84);
not(t_3819, k6);
and(x85, t_3818, t_3819);
not(t_3820, f85);
not(t_3821, x8);
and(y85, t_3820, t_3821);
not(t_3822, w84);
not(t_3823, n9);
and(z85, t_3822, t_3823);
not(t_3824, z84);
not(t_3825, c84);
and(a86, t_3824, t_3825);
not(t_3826, a85);
not(t_3827, e84);
and(b86, t_3826, t_3827);
not(t_3828, b85);
not(t_3829, g84);
and(c86, t_3828, t_3829);
not(t_3830, h85);
not(t_3831, i85);
and(d86, t_3830, t_3831);
not(t_3832, m84);
not(t_3833, j85);
and(e86, t_3832, t_3833);
not(t_3834, j85);
not(t_3835, n84);
and(f86, t_3834, t_3835);
not(t_3836, k85);
not(t_3837, l85);
and(g86, t_3836, t_3837);
not(t_3838, m85);
not(t_3839, w85);
and(h86, t_3838, t_3839);
not(t_3840, k82);
not(t_3841, x85);
and(i86, t_3840, t_3841);
not(t_3842, p84);
not(t_3843, x85);
and(j86, t_3842, t_3843);
not(t_3844, o85);
not(t_3845, p85);
and(k86, t_3844, t_3845);
not(t_3846, t84);
not(t_3847, q85);
and(l86, t_3846, t_3847);
not(t_3848, q85);
not(t_3849, u84);
and(m86, t_3848, t_3849);
not(t_3850, r85);
not(t_3851, s85);
and(n86, t_3850, t_3851);
not(t_3852, t85);
not(t_3853, y85);
and(o86, t_3852, t_3853);
not(t_3854, r82);
not(t_3855, z85);
and(p86, t_3854, t_3855);
not(t_3856, w84);
not(t_3857, z85);
and(q86, t_3856, t_3857);
not(t_3858, v85);
not(t_3859, a86);
and(r86, t_3858, t_3859);
not(t_3860, a85);
not(t_3861, b86);
and(s86, t_3860, t_3861);
not(t_3862, b85);
not(t_3863, c86);
and(t86, t_3862, t_3863);
not(t_3864, x85);
not(t_3865, k6);
and(u86, t_3864, t_3865);
not(t_3866, n85);
not(t_3867, a7);
and(v86, t_3866, t_3867);
not(t_3868, z85);
not(t_3869, n9);
and(w86, t_3868, t_3869);
not(t_3870, u85);
not(t_3871, d10);
and(x86, t_3870, t_3871);
not(t_3872, b86);
not(t_3873, e84);
and(y86, t_3872, t_3873);
not(t_3874, c86);
not(t_3875, g84);
and(z86, t_3874, t_3875);
not(t_3876, e86);
not(t_3877, f86);
and(a87, t_3876, t_3877);
not(t_3878, k85);
not(t_3879, g86);
and(b87, t_3878, t_3879);
not(t_3880, g86);
not(t_3881, l85);
and(c87, t_3880, t_3881);
not(t_3882, h86);
not(t_3883, i86);
and(d87, t_3882, t_3883);
not(t_3884, j86);
not(t_3885, u86);
and(e87, t_3884, t_3885);
not(t_3886, m83);
not(t_3887, v86);
and(f87, t_3886, t_3887);
not(t_3888, n85);
not(t_3889, v86);
and(g87, t_3888, t_3889);
not(t_3890, l86);
not(t_3891, m86);
and(h87, t_3890, t_3891);
not(t_3892, r85);
not(t_3893, n86);
and(i87, t_3892, t_3893);
not(t_3894, n86);
not(t_3895, s85);
and(j87, t_3894, t_3895);
not(t_3896, o86);
not(t_3897, p86);
and(k87, t_3896, t_3897);
not(t_3898, q86);
not(t_3899, w86);
and(l87, t_3898, t_3899);
not(t_3900, t83);
not(t_3901, x86);
and(m87, t_3900, t_3901);
not(t_3902, u85);
not(t_3903, x86);
and(n87, t_3902, t_3903);
not(t_3904, s86);
not(t_3905, y86);
and(o87, t_3904, t_3905);
not(t_3906, t86);
not(t_3907, z86);
and(p87, t_3906, t_3907);
not(t_3908, v86);
not(t_3909, a7);
and(q87, t_3908, t_3909);
not(t_3910, k86);
not(t_3911, q7);
and(r87, t_3910, t_3911);
not(t_3912, x86);
not(t_3913, d10);
and(s87, t_3912, t_3913);
not(t_3914, r86);
not(t_3915, t10);
and(t87, t_3914, t_3915);
not(t_3916, b87);
not(t_3917, c87);
and(u87, t_3916, t_3917);
not(t_3918, h86);
not(t_3919, d87);
and(v87, t_3918, t_3919);
not(t_3920, d87);
not(t_3921, i86);
and(w87, t_3920, t_3921);
not(t_3922, e87);
not(t_3923, f87);
and(x87, t_3922, t_3923);
not(t_3924, g87);
not(t_3925, q87);
and(y87, t_3924, t_3925);
not(t_3926, s84);
not(t_3927, r87);
and(z87, t_3926, t_3927);
not(t_3928, k86);
not(t_3929, r87);
and(a88, t_3928, t_3929);
not(t_3930, i87);
not(t_3931, j87);
and(b88, t_3930, t_3931);
not(t_3932, o86);
not(t_3933, k87);
and(c88, t_3932, t_3933);
not(t_3934, k87);
not(t_3935, p86);
and(d88, t_3934, t_3935);
not(t_3936, l87);
not(t_3937, m87);
and(e88, t_3936, t_3937);
not(t_3938, n87);
not(t_3939, s87);
and(f88, t_3938, t_3939);
not(t_3940, z84);
not(t_3941, t87);
and(g88, t_3940, t_3941);
not(t_3942, r86);
not(t_3943, t87);
and(h88, t_3942, t_3943);
not(t_3944, r87);
not(t_3945, q7);
and(i88, t_3944, t_3945);
not(t_3946, h87);
not(t_3947, g8);
and(j88, t_3946, t_3947);
not(t_3948, t87);
not(t_3949, t10);
and(k88, t_3948, t_3949);
not(t_3950, o87);
not(t_3951, j11);
and(l88, t_3950, t_3951);
not(t_3952, p87);
not(t_3953, z11);
and(m88, t_3952, t_3953);
not(t_3954, v87);
not(t_3955, w87);
and(n88, t_3954, t_3955);
not(t_3956, e87);
not(t_3957, x87);
and(o88, t_3956, t_3957);
not(t_3958, x87);
not(t_3959, f87);
and(p88, t_3958, t_3959);
not(t_3960, y87);
not(t_3961, z87);
and(q88, t_3960, t_3961);
not(t_3962, a88);
not(t_3963, i88);
and(r88, t_3962, t_3963);
not(t_3964, q85);
not(t_3965, j88);
and(s88, t_3964, t_3965);
not(t_3966, h87);
not(t_3967, j88);
and(t88, t_3966, t_3967);
not(t_3968, c88);
not(t_3969, d88);
and(u88, t_3968, t_3969);
not(t_3970, l87);
not(t_3971, e88);
and(v88, t_3970, t_3971);
not(t_3972, e88);
not(t_3973, m87);
and(w88, t_3972, t_3973);
not(t_3974, f88);
not(t_3975, g88);
and(x88, t_3974, t_3975);
not(t_3976, h88);
not(t_3977, k88);
and(y88, t_3976, t_3977);
not(t_3978, o87);
not(t_3979, l88);
and(z88, t_3978, t_3979);
not(t_3980, p87);
not(t_3981, m88);
and(a89, t_3980, t_3981);
not(t_3982, j88);
not(t_3983, g8);
and(b89, t_3982, t_3983);
not(t_3984, b88);
not(t_3985, w8);
and(c89, t_3984, t_3985);
not(t_3986, b86);
not(t_3987, l88);
and(d89, t_3986, t_3987);
not(t_3988, l88);
not(t_3989, j11);
and(e89, t_3988, t_3989);
not(t_3990, c86);
not(t_3991, m88);
and(f89, t_3990, t_3991);
not(t_3992, m88);
not(t_3993, z11);
and(g89, t_3992, t_3993);
not(t_3994, o88);
not(t_3995, p88);
and(h89, t_3994, t_3995);
not(t_3996, y87);
not(t_3997, q88);
and(i89, t_3996, t_3997);
not(t_3998, q88);
not(t_3999, z87);
and(j89, t_3998, t_3999);
not(t_4000, r88);
not(t_4001, s88);
and(k89, t_4000, t_4001);
not(t_4002, t88);
not(t_4003, b89);
and(l89, t_4002, t_4003);
not(t_4004, n86);
not(t_4005, c89);
and(m89, t_4004, t_4005);
not(t_4006, b88);
not(t_4007, c89);
and(n89, t_4006, t_4007);
not(t_4008, v88);
not(t_4009, w88);
and(o89, t_4008, t_4009);
not(t_4010, f88);
not(t_4011, x88);
and(p89, t_4010, t_4011);
not(t_4012, x88);
not(t_4013, g88);
and(q89, t_4012, t_4013);
not(t_4014, y88);
not(t_4015, d89);
and(r89, t_4014, t_4015);
not(t_4016, z88);
not(t_4017, e89);
and(s89, t_4016, t_4017);
not(t_4018, c89);
not(t_4019, w8);
and(t89, t_4018, t_4019);
not(t_4020, u88);
not(t_4021, m9);
and(u89, t_4020, t_4021);
not(t_4022, i89);
not(t_4023, j89);
and(v89, t_4022, t_4023);
not(t_4024, r88);
not(t_4025, k89);
and(w89, t_4024, t_4025);
not(t_4026, k89);
not(t_4027, s88);
and(x89, t_4026, t_4027);
not(t_4028, l89);
not(t_4029, m89);
and(y89, t_4028, t_4029);
not(t_4030, n89);
not(t_4031, t89);
and(z89, t_4030, t_4031);
not(t_4032, k87);
not(t_4033, u89);
and(a90, t_4032, t_4033);
not(t_4034, u88);
not(t_4035, u89);
and(b90, t_4034, t_4035);
not(t_4036, p89);
not(t_4037, q89);
and(c90, t_4036, t_4037);
not(t_4038, y88);
not(t_4039, r89);
and(d90, t_4038, t_4039);
not(t_4040, u89);
not(t_4041, m9);
and(e90, t_4040, t_4041);
not(t_4042, o89);
not(t_4043, c10);
and(f90, t_4042, t_4043);
not(t_4044, r89);
not(t_4045, d89);
and(g90, t_4044, t_4045);
not(t_4046, s89);
not(t_4047, f89);
and(h90, t_4046, t_4047);
not(t_4048, w89);
not(t_4049, x89);
and(i90, t_4048, t_4049);
not(t_4050, l89);
not(t_4051, y89);
and(j90, t_4050, t_4051);
not(t_4052, y89);
not(t_4053, m89);
and(k90, t_4052, t_4053);
not(t_4054, z89);
not(t_4055, a90);
and(l90, t_4054, t_4055);
not(t_4056, b90);
not(t_4057, e90);
and(m90, t_4056, t_4057);
not(t_4058, e88);
not(t_4059, f90);
and(n90, t_4058, t_4059);
not(t_4060, o89);
not(t_4061, f90);
and(o90, t_4060, t_4061);
not(t_4062, d90);
not(t_4063, g90);
and(p90, t_4062, t_4063);
not(t_4064, s89);
not(t_4065, h90);
and(q90, t_4064, t_4065);
not(t_4066, f90);
not(t_4067, c10);
and(r90, t_4066, t_4067);
not(t_4068, c90);
not(t_4069, s10);
and(s90, t_4068, t_4069);
not(t_4070, h90);
not(t_4071, f89);
and(t90, t_4070, t_4071);
not(t_4072, j90);
not(t_4073, k90);
and(u90, t_4072, t_4073);
not(t_4074, z89);
not(t_4075, l90);
and(v90, t_4074, t_4075);
not(t_4076, l90);
not(t_4077, a90);
and(w90, t_4076, t_4077);
not(t_4078, m90);
not(t_4079, n90);
and(x90, t_4078, t_4079);
not(t_4080, o90);
not(t_4081, r90);
and(y90, t_4080, t_4081);
not(t_4082, x88);
not(t_4083, s90);
and(z90, t_4082, t_4083);
not(t_4084, c90);
not(t_4085, s90);
and(a91, t_4084, t_4085);
not(t_4086, q90);
not(t_4087, t90);
and(b91, t_4086, t_4087);
not(t_4088, s90);
not(t_4089, s10);
and(c91, t_4088, t_4089);
not(t_4090, p90);
not(t_4091, i11);
and(d91, t_4090, t_4091);
not(t_4092, v90);
not(t_4093, w90);
and(e91, t_4092, t_4093);
not(t_4094, m90);
not(t_4095, x90);
and(f91, t_4094, t_4095);
not(t_4096, x90);
not(t_4097, n90);
and(g91, t_4096, t_4097);
not(t_4098, y90);
not(t_4099, z90);
and(h91, t_4098, t_4099);
not(t_4100, a91);
not(t_4101, c91);
and(i91, t_4100, t_4101);
not(t_4102, r89);
not(t_4103, d91);
and(j91, t_4102, t_4103);
not(t_4104, p90);
not(t_4105, d91);
and(k91, t_4104, t_4105);
not(t_4106, d91);
not(t_4107, i11);
and(l91, t_4106, t_4107);
not(t_4108, b91);
not(t_4109, y11);
and(m91, t_4108, t_4109);
not(t_4110, f91);
not(t_4111, g91);
and(n91, t_4110, t_4111);
not(t_4112, y90);
not(t_4113, h91);
and(o91, t_4112, t_4113);
not(t_4114, h91);
not(t_4115, z90);
and(p91, t_4114, t_4115);
not(t_4116, i91);
not(t_4117, j91);
and(q91, t_4116, t_4117);
not(t_4118, k91);
not(t_4119, l91);
and(r91, t_4118, t_4119);
not(t_4120, b91);
not(t_4121, m91);
and(s91, t_4120, t_4121);
not(t_4122, h90);
not(t_4123, m91);
and(t91, t_4122, t_4123);
not(t_4124, m91);
not(t_4125, y11);
and(u91, t_4124, t_4125);
not(t_4126, o91);
not(t_4127, p91);
and(v91, t_4126, t_4127);
not(t_4128, i91);
not(t_4129, q91);
and(w91, t_4128, t_4129);
not(t_4130, q91);
not(t_4131, j91);
and(x91, t_4130, t_4131);
not(t_4132, r91);
not(t_4133, t91);
and(y91, t_4132, t_4133);
not(t_4134, w91);
not(t_4135, x91);
and(z91, t_4134, t_4135);
not(t_4136, r91);
not(t_4137, y91);
and(a92, t_4136, t_4137);
not(t_4138, y91);
not(t_4139, t91);
and(b92, t_4138, t_4139);
not(t_4140, a92);
not(t_4141, b92);
and(c92, t_4140, t_4141);
not(d92, c92);
not(t_4142, y91);
not(t_4143, d92);
and(e92, t_4142, t_4143);
not(t_4144, c92);
not(t_4145, d92);
and(f92, t_4144, t_4145);
not(g92, d92);
not(t_4146, z91);
not(t_4147, e92);
and(h92, t_4146, t_4147);
not(t_4148, q91);
not(t_4149, h92);
and(i92, t_4148, t_4149);
not(t_4150, z91);
not(t_4151, h92);
and(j92, t_4150, t_4151);
not(t_4152, h92);
not(t_4153, e92);
and(k92, t_4152, t_4153);
not(t_4154, v91);
not(t_4155, i92);
and(l92, t_4154, t_4155);
not(t_4156, h91);
not(t_4157, l92);
and(m92, t_4156, t_4157);
not(t_4158, v91);
not(t_4159, l92);
and(n92, t_4158, t_4159);
not(t_4160, l92);
not(t_4161, i92);
and(o92, t_4160, t_4161);
not(t_4162, n91);
not(t_4163, m92);
and(p92, t_4162, t_4163);
not(t_4164, x90);
not(t_4165, p92);
and(q92, t_4164, t_4165);
not(t_4166, n91);
not(t_4167, p92);
and(r92, t_4166, t_4167);
not(t_4168, p92);
not(t_4169, m92);
and(s92, t_4168, t_4169);
not(t_4170, e91);
not(t_4171, q92);
and(t92, t_4170, t_4171);
not(t_4172, l90);
not(t_4173, t92);
and(u92, t_4172, t_4173);
not(t_4174, e91);
not(t_4175, t92);
and(v92, t_4174, t_4175);
not(t_4176, t92);
not(t_4177, q92);
and(w92, t_4176, t_4177);
not(t_4178, u90);
not(t_4179, u92);
and(x92, t_4178, t_4179);
not(t_4180, y89);
not(t_4181, x92);
and(y92, t_4180, t_4181);
not(t_4182, u90);
not(t_4183, x92);
and(z92, t_4182, t_4183);
not(t_4184, x92);
not(t_4185, u92);
and(a93, t_4184, t_4185);
not(t_4186, i90);
not(t_4187, y92);
and(b93, t_4186, t_4187);
not(t_4188, k89);
not(t_4189, b93);
and(c93, t_4188, t_4189);
not(t_4190, i90);
not(t_4191, b93);
and(d93, t_4190, t_4191);
not(t_4192, b93);
not(t_4193, y92);
and(e93, t_4192, t_4193);
not(t_4194, v89);
not(t_4195, c93);
and(f93, t_4194, t_4195);
not(t_4196, q88);
not(t_4197, f93);
and(g93, t_4196, t_4197);
not(t_4198, v89);
not(t_4199, f93);
and(h93, t_4198, t_4199);
not(t_4200, f93);
not(t_4201, c93);
and(i93, t_4200, t_4201);
not(t_4202, h89);
not(t_4203, g93);
and(j93, t_4202, t_4203);
not(t_4204, x87);
not(t_4205, j93);
and(k93, t_4204, t_4205);
not(t_4206, h89);
not(t_4207, j93);
and(l93, t_4206, t_4207);
not(t_4208, j93);
not(t_4209, g93);
and(m93, t_4208, t_4209);
not(t_4210, n88);
not(t_4211, k93);
and(n93, t_4210, t_4211);
not(t_4212, d87);
not(t_4213, n93);
and(o93, t_4212, t_4213);
not(t_4214, n88);
not(t_4215, n93);
and(p93, t_4214, t_4215);
not(t_4216, n93);
not(t_4217, k93);
and(q93, t_4216, t_4217);
not(t_4218, u87);
not(t_4219, o93);
and(r93, t_4218, t_4219);
not(t_4220, g86);
not(t_4221, r93);
and(s93, t_4220, t_4221);
not(t_4222, u87);
not(t_4223, r93);
and(t93, t_4222, t_4223);
not(t_4224, r93);
not(t_4225, o93);
and(u93, t_4224, t_4225);
not(t_4226, a87);
not(t_4227, s93);
and(v93, t_4226, t_4227);
not(t_4228, j85);
not(t_4229, v93);
and(w93, t_4228, t_4229);
not(t_4230, a87);
not(t_4231, v93);
and(x93, t_4230, t_4231);
not(t_4232, v93);
not(t_4233, s93);
and(y93, t_4232, t_4233);
not(t_4234, d86);
not(t_4235, w93);
and(z93, t_4234, t_4235);
not(t_4236, l84);
not(t_4237, z93);
and(a94, t_4236, t_4237);
not(t_4238, d86);
not(t_4239, z93);
and(b94, t_4238, t_4239);
not(t_4240, z93);
not(t_4241, w93);
and(c94, t_4240, t_4241);
not(t_4242, g85);
not(t_4243, a94);
and(d94, t_4242, t_4243);
not(t_4244, f83);
not(t_4245, d94);
and(e94, t_4244, t_4245);
not(t_4246, g85);
not(t_4247, d94);
and(f94, t_4246, t_4247);
not(t_4248, d94);
not(t_4249, a94);
and(g94, t_4248, t_4249);
not(t_4250, i84);
not(t_4251, e94);
and(h94, t_4250, t_4251);
not(t_4252, i84);
not(t_4253, h94);
and(i94, t_4252, t_4253);
not(t_4254, h94);
not(t_4255, e94);
and(j94, t_4254, t_4255);
endmodule
module top;
	parameter in_width = 32,
		patterns = 5000,
		step = 1;
	reg [1:in_width] in_mem[1:patterns];
	integer index;

	wire i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,
		i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,
		i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,
		i30,i31;

	assign {i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,
		i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,
		i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,
		i30,i31} = 
		$getpattern(in_mem[index]);

	initial $monitor($time,,o0,o1,o2,o3,o4,o5,o6,o7,o8,o9,
		o10,o11,o12,o13,o14,o15,o16,o17,o18,o19,
		o20,o21,o22,o23,o24,o25,o26,o27,o28,o29,
		o30,o31);
	initial
		begin
			$readmemb("patt.mem", in_mem);
			for(index = 1; index <= patterns; index = index + 1)
				#step;
		end

	foobar cct(o0,o1,o2,o3,o4,o5,o6,o7,o8,o9,
		o10,o11,o12,o13,o14,o15,o16,o17,o18,o19,
		o20,o21,o22,o23,o24,o25,o26,o27,o28,o29,
		o30,o31,i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,
		i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,
		i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,
		i30,i31);
endmodule
