// IWLS benchmark module "CM162" printed on Wed May 29 16:07:20 2002
module CM162(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s);
input
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n;
output
  o,
  p,
  q,
  r,
  s;
wire
  \[7] ,
  p0,
  e0,
  q0,
  f0,
  r0,
  \[0] ,
  \[11] ,
  \[1] ,
  \[2] ,
  \[13] ,
  \[3] ,
  \[4] ,
  \[5] ;
assign
  \[7]  = (e0 & k) | ((k & i) | (r0 | ~f0)),
  p0 = (~l & ~r0) | (l & r0),
  e0 = (~\[11]  & i) | (\[11]  & ~i),
  q0 = (~\[13]  & m) | (\[13]  & ~m),
  f0 = (~\[4]  & (f & d)) | (f & (d & ~c)),
  r0 = ~\[11]  & (~k & ~i),
  \[0]  = (\[5]  & ~f0) | ((\[5]  & ~e0) | ((~f0 & ~a) | (~e0 & ~a))),
  \[11]  = ~e | (~d | ~c),
  \[1]  = (\[7]  & \[5] ) | (\[7]  & ~b),
  o = \[0] ,
  p = \[1] ,
  q = \[2] ,
  r = \[3] ,
  s = \[4] ,
  \[2]  = (\[5]  & ~p0) | ((\[5]  & ~f0) | ((~p0 & ~g) | (~f0 & ~g))),
  \[13]  = ~r0 | l,
  \[3]  = (\[5]  & ~q0) | ((\[5]  & ~f0) | ((~q0 & ~h) | (~f0 & ~h))),
  \[4]  = n & (j & e),
  \[5]  = ~f | d;
endmodule

