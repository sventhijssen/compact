// IWLS benchmark module "term1" printed on Wed May 29 16:09:31 2002
module term1(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, \x , y, z, a0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0);
input
  g0,
  h0,
  i0,
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  t,
  u,
  v,
  w,
  \x ,
  y,
  z,
  a0,
  c0,
  d0,
  e0,
  f0;
output
  j0,
  k0,
  l0,
  m0,
  n0,
  o0,
  p0,
  q0,
  r0,
  s0;
wire
  f5,
  \[26] ,
  \[27] ,
  i7,
  \[43] ,
  \[10] ,
  \[45] ,
  \[11] ,
  \[46] ,
  \[12] ,
  n4,
  \[48] ,
  \[14] ,
  p4,
  \[0] ,
  \[15] ,
  \[30] ,
  \[1] ,
  \[2] ,
  \[17] ,
  \[3] ,
  s5,
  \[18] ,
  \[33] ,
  \[4] ,
  \[5] ,
  \[6] ,
  \[7] ,
  w5,
  \[8] ,
  \[9] ,
  z2,
  \[39] ,
  \[21] ,
  b7,
  c3,
  \[22] ,
  c6,
  \[23] ;
assign
  f5 = ~c0 & ~d0,
  \[26]  = \[21]  | ~d,
  \[27]  = ~g | c,
  i7 = (~\[48]  & ~b7) | ((\[48]  & b7) | ~\[26] ),
  \[43]  = (~\[18]  & (n4 & r)) | ((\[23]  & ~r) | ((\[22]  & ~q) | ((\[18]  & ~s5) | ~\[12] ))),
  j0 = \[0] ,
  k0 = \[1] ,
  \[10]  = ~a0 & a,
  \[45]  = z2 | ~f0,
  l0 = \[2] ,
  \[11]  = (~w & ~r) | ((~v & ~q) | (~u & ~p)),
  \[46]  = p4 | ~g0,
  m0 = \[3] ,
  \[12]  = t | s,
  n0 = \[4] ,
  n4 = (t & ~n) | ((s & ~o) | w5),
  \[48]  = f | d,
  o0 = \[5] ,
  \[14]  = ~d | ~c,
  p0 = \[6] ,
  p4 = (~\[39]  & f0) | (\[39]  & ~f0),
  \[0]  = ~h0,
  \[15]  = (\[18]  & (s5 & (q & k))) | ((~\[23]  & (~\[18]  & ~s5)) | (~\[22]  & (\[18]  & s5))),
  q0 = \[7] ,
  \[30]  = (~\[11]  & c3) | (\[17]  | ~\[14] ),
  \[1]  = (~i0 & (~d & ~c)) | ((~h0 & (~d & c)) | ((~h0 & (d & ~c)) | (~\[14]  & ~i0))),
  r0 = \[8] ,
  \[2]  = (\[26]  & (~b7 & (~j & (i & (~c & b))))) | ((~\[27]  & (i7 & (~j & (i & ~b)))) | ((\[27]  & (~i7 & (~j & (i & ~b)))) | ((~\[21]  & (~\[14]  & (~j & (i & b)))) | (b7 & (~j & (i & (c & b))))))),
  \[17]  = a0 | (~z | ~b),
  s0 = \[9] ,
  \[3]  = ~\[30]  & ~c0,
  s5 = w5 & r,
  \[18]  = ~q | ~p,
  \[33]  = y | t,
  \[4]  = (~\[30]  & (~f5 & ~d0)) | (~f5 & \[3] ),
  \[5]  = (~\[30]  & (z2 & (~\[4]  & ~\[3] ))) | (~\[30]  & (z2 & e0)),
  \[6]  = (~\[30]  & (~z2 & ~f0)) | (~\[30]  & (z2 & f0)),
  \[7]  = (~\[45]  & ~g0) | ((\[45]  & g0) | \[30] ),
  w5 = s & t,
  \[8]  = (~\[46]  & (~\[43]  & (~\[18]  & (\[10]  & ~h0)))) | ((~\[46]  & (\[15]  & (\[10]  & ~h0))) | ((~\[15]  & (\[10]  & (h0 & ~p))) | ((\[46]  & (\[10]  & h0)) | (\[43]  & (\[10]  & h0))))),
  \[9]  = (~\[43]  & (~\[39]  & (\[10]  & (~i0 & (g0 & (f0 & p)))))) | ((~\[43]  & (\[39]  & (\[10]  & (p4 & (~i0 & (~g0 & p)))))) | ((~\[39]  & (\[15]  & (\[10]  & (~i0 & (g0 & f0))))) | ((\[39]  & (\[15]  & (\[10]  & (p4 & (~i0 & ~g0))))) | ((~\[39]  & (\[10]  & (i0 & ~g0))) | ((\[18]  & (~\[15]  & (\[10]  & i0))) | ((\[10]  & (i0 & (g0 & ~f0))) | ((\[43]  & (\[10]  & i0)) | (\[10]  & (~p4 & i0))))))))),
  z2 = ~c0 | (~d0 | ~e0),
  \[39]  = f5 | ~e0,
  \[21]  = ~h | ~e,
  b7 = (~h & (~e & d)) | ((~h & (e & ~d)) | (h & (~e & ~d))),
  c3 = (\[33]  & \x ) | (\[33]  & s),
  \[22]  = ~p | ~l,
  c6 = 0,
  \[23]  = ~w5 | ~m;
endmodule

