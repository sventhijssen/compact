// IWLS benchmark module "pm1" printed on Wed May 29 16:09:22 2002
module pm1(a, b, c, d, e, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, \x , y, z, a0, b0, c0, d0);
input
  a,
  b,
  c,
  d,
  e,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q;
output
  c0,
  d0,
  r,
  s,
  t,
  u,
  v,
  w,
  \x ,
  y,
  z,
  a0,
  b0;
wire
  \[7] ,
  \[18] ,
  \[8] ,
  \[9] ,
  \[10] ,
  \[0] ,
  \[11] ,
  \[1] ,
  \[12] ,
  \[2] ,
  \[3] ,
  \[14] ,
  \[4] ,
  \[15] ,
  \[5] ,
  \[6] ,
  \[17] ;
assign
  c0 = \[11] ,
  \[7]  = ~q,
  \[18]  = \[9]  & n,
  d0 = \[12] ,
  \[8]  = (~\[12]  & (~\[10]  & \[9] )) | \[17] ,
  \[9]  = (~\[15]  & (~n & ~m)) | (~\[17]  & n),
  \[10]  = \[18]  & (\[14]  & ~\[12] ),
  \[0]  = b | (m | n),
  \[11]  = (~\[17]  & (~\[9]  & ~b)) | (\[18]  & \[6] ),
  \[1]  = m | ~n,
  \[12]  = \[18]  & ~k,
  r = \[0] ,
  s = \[1] ,
  t = \[2] ,
  \[2]  = ~n | (~m | (~k | (~j | (~i | (~h | ~g))))),
  u = \[3] ,
  v = \[4] ,
  w = \[5] ,
  \x  = \[6] ,
  y = \[7] ,
  z = \[8] ,
  \[3]  = ~\[2]  | (~\[1]  | (~n | ~k)),
  \[14]  = ~e | (~d | ~c),
  \[4]  = ~p,
  \[15]  = l | ~a,
  a0 = \[9] ,
  \[5]  = ~o,
  b0 = \[10] ,
  \[6]  = (\[14]  & (k & b)) | (~\[1]  & (k & b)),
  \[17]  = \[15]  | ~m;
endmodule

