module foobar(h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x, y, z, a0, b0, c0, d0, e0, f0, g0);
input a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x, y, z, a0, b0, c0, d0, e0, f0, g0;
output h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1;
not(t_0, e33);
not(t_1, k32);
or(h0, t_0, t_1);
not(t_2, d33);
not(t_3, j32);
or(i0, t_2, t_3);
not(t_4, c33);
not(t_5, i32);
or(j0, t_4, t_5);
not(t_6, b33);
not(t_7, h32);
or(k0, t_6, t_7);
not(t_8, v32);
not(t_9, b32);
or(l0, t_8, t_9);
not(t_10, q32);
not(t_11, w31);
or(m0, t_10, t_11);
not(t_12, p32);
not(t_13, v31);
or(n0, t_12, t_13);
not(t_14, a33);
not(t_15, g32);
or(o0, t_14, t_15);
not(t_16, z32);
not(t_17, f32);
or(p0, t_16, t_17);
not(t_18, y32);
not(t_19, e32);
or(q0, t_18, t_19);
not(t_20, x32);
not(t_21, d32);
or(r0, t_20, t_21);
not(t_22, w32);
not(t_23, c32);
or(s0, t_22, t_23);
not(t_24, u32);
not(t_25, a32);
or(t0, t_24, t_25);
not(t_26, t32);
not(t_27, z31);
or(u0, t_26, t_27);
not(t_28, s32);
not(t_29, y31);
or(v0, t_28, t_29);
not(t_30, r32);
not(t_31, x31);
or(w0, t_30, t_31);
not(t_32, l29);
not(t_33, j33);
and(x0, t_32, t_33);
and(y0, r34, l4);
and(z0, m4, q34);
and(a1, o4, v34);
and(b1, t34, p4);
and(c1, q4, s34);
not(t_34, w34);
not(t_35, o34);
or(d1, t_34, t_35);
not(t_36, x34);
not(t_37, p34);
or(e1, t_36, t_37);
and(f1, b35, n4);
not(f2, g0);
buf(g2, g0);
buf(h2, g0);
not(i2, g0);
buf(j2, g0);
not(k2, g0);
not(l2, g0);
not(m2, f0);
not(n2, f0);
buf(o2, f0);
not(p2, e0);
buf(q2, e0);
not(r2, e0);
buf(s2, e0);
not(t2, d0);
not(u2, c0);
not(v2, b0);
not(w2, a0);
not(x2, z);
not(y2, y);
not(z2, x);
not(a3, x);
buf(b3, w);
buf(c3, w);
not(t_38, d0);
not(t_39, v);
or(d3, t_38, t_39);
not(t_40, c0);
not(t_41, u);
or(e3, t_40, t_41);
not(f3, p);
buf(g3, p);
not(h3, o);
buf(i3, o);
not(j3, n);
buf(k3, n);
not(l3, m);
buf(m3, m);
not(n3, l);
buf(o3, l);
not(p3, k);
buf(q3, k);
not(r3, j);
buf(s3, j);
not(t3, i);
buf(u3, i);
not(v3, h);
buf(w3, h);
not(x3, g);
buf(y3, g);
not(z3, f);
buf(a4, f);
not(b4, e);
buf(c4, e);
not(d4, d);
buf(e4, d);
not(f4, c);
buf(g4, c);
not(h4, b);
buf(i4, b);
not(j4, a);
buf(k4, a);
not(t_42, g2);
not(t_43, n2);
or(l4, t_42, t_43);
not(t_44, g2);
not(t_45, n2);
or(m4, t_44, t_45);
not(t_46, g2);
not(t_47, n2);
or(n4, t_46, t_47);
not(t_48, g2);
not(t_49, n2);
or(o4, t_48, t_49);
not(t_50, g2);
not(t_51, n2);
or(p4, t_50, t_51);
not(t_52, g2);
not(t_53, n2);
or(q4, t_52, t_53);
not(t_54, u2);
not(t_55, h2);
or(r4, t_54, t_55);
not(t_56, t2);
not(t_57, h2);
or(s4, t_56, t_57);
and(t4, e3, j2);
and(u4, d3, j2);
not(t_58, p2);
not(t_59, b3);
or(v4, t_58, t_59);
not(t_60, p2);
not(t_61, z2);
or(w4, t_60, t_61);
buf(x4, v2);
buf(y4, v2);
buf(z4, w2);
buf(a5, w2);
buf(b5, x2);
buf(c5, x2);
buf(d5, y2);
buf(e5, y2);
not(t_62, x);
not(t_63, b3);
or(f5, t_62, t_63);
and(g5, v, i2);
and(h5, u, i2);
and(i5, t, c3, i2);
and(j5, s, c3, i2);
and(k5, r, a3, i2);
and(l5, q, a3, i2);
buf(m5, f3);
buf(n5, f3);
buf(o5, f3);
not(p5, g3);
buf(q5, h3);
buf(r5, h3);
buf(s5, h3);
not(t5, i3);
buf(u5, j3);
buf(v5, j3);
buf(w5, j3);
not(x5, k3);
buf(y5, l3);
buf(z5, l3);
buf(a6, l3);
not(b6, m3);
buf(c6, n3);
buf(d6, n3);
not(e6, o3);
buf(f6, p3);
buf(g6, p3);
not(h6, q3);
buf(i6, r3);
buf(j6, r3);
buf(k6, r3);
not(l6, s3);
buf(m6, t3);
buf(n6, t3);
buf(o6, t3);
buf(p6, t3);
not(q6, u3);
buf(r6, v3);
buf(s6, v3);
buf(t6, v3);
not(u6, w3);
buf(v6, x3);
buf(w6, x3);
buf(x6, x3);
not(y6, y3);
buf(z6, z3);
buf(a7, z3);
not(b7, a4);
buf(c7, b4);
buf(d7, b4);
not(e7, c4);
buf(f7, d4);
buf(g7, d4);
buf(h7, d4);
buf(i7, d4);
not(j7, e4);
buf(k7, f4);
buf(l7, f4);
buf(m7, f4);
not(n7, g4);
buf(o7, h4);
buf(p7, h4);
not(q7, i4);
buf(r7, j4);
buf(s7, j4);
buf(t7, j4);
not(u7, k4);
and(v7, o2, f2, f5);
not(t_64, f5);
not(t_65, f2);
not(t_66, o2);
or(w7, t_64, t_65, t_66);
not(t_67, f5);
not(t_68, h2);
not(t_69, q2);
not(t_70, u2);
or(x7, t_67, t_68, t_69, t_70);
not(t_71, f5);
not(t_72, h2);
not(t_73, q2);
not(t_74, t2);
or(y7, t_71, t_72, t_73, t_74);
not(z7, t4);
not(a8, u4);
not(b8, x4);
not(c8, y4);
not(d8, z4);
not(e8, a5);
not(f8, b5);
not(g8, c5);
not(h8, d5);
not(i8, e5);
buf(j8, g5);
buf(k8, g5);
buf(l8, h5);
buf(m8, h5);
not(t_75, v4);
not(t_76, t);
or(n8, t_75, t_76);
not(o8, i5);
not(t_77, v4);
not(t_78, s);
or(p8, t_77, t_78);
and(q8, s, v4);
not(r8, j5);
not(t_79, w4);
not(t_80, r);
or(s8, t_79, t_80);
not(t8, k5);
not(t_81, w4);
not(t_82, q);
or(u8, t_81, t_82);
and(v8, q, w4);
buf(w8, l5);
buf(x8, l5);
not(y8, m5);
not(z8, n5);
buf(a9, o5);
buf(b9, o5);
buf(c9, q5);
buf(d9, q5);
not(e9, r5);
not(f9, s5);
buf(g9, u5);
buf(h9, u5);
not(i9, v5);
buf(j9, w5);
buf(k9, w5);
not(l9, y5);
not(m9, z5);
not(n9, a6);
buf(o9, c6);
buf(p9, c6);
not(q9, d6);
buf(r9, f6);
buf(s9, f6);
not(t9, g6);
buf(u9, i6);
buf(v9, i6);
not(w9, j6);
not(x9, k6);
buf(y9, m6);
buf(z9, m6);
not(a10, n6);
not(b10, o6);
not(c10, p6);
not(d10, r6);
not(e10, s6);
not(f10, t6);
not(g10, v6);
not(h10, w6);
not(i10, x6);
buf(j10, z6);
buf(k10, z6);
not(l10, a7);
buf(m10, c7);
buf(n10, c7);
not(o10, d7);
not(p10, f7);
not(q10, g7);
not(r10, h7);
not(s10, i7);
not(t10, k7);
not(u10, l7);
not(v10, m7);
buf(w10, o7);
buf(x10, o7);
not(y10, p7);
buf(z10, r7);
buf(a11, r7);
not(b11, s7);
not(c11, t7);
not(t_83, w7);
not(t_84, x7);
or(d11, t_83, t_84);
not(t_85, w7);
not(t_86, y7);
or(e11, t_85, t_86);
not(f11, j8);
not(g11, k8);
not(h11, l8);
not(i11, m8);
not(j11, n8);
buf(k11, n8);
not(t_87, n9);
not(t_88, i5);
or(l11, t_87, t_88);
buf(m11, p8);
buf(n11, p8);
not(o11, s8);
buf(p11, s8);
not(t_89, e9);
not(t_90, k5);
or(q11, t_89, t_90);
buf(r11, u8);
buf(s11, u8);
not(t11, w8);
not(t_91, b11);
not(t_92, w8);
or(u11, t_91, t_92);
not(t_93, c11);
not(t_94, x8);
or(v11, t_93, t_94);
not(w11, x8);
not(t_95, y8);
not(t_96, c9);
or(x11, t_95, t_96);
not(t_97, z8);
not(t_98, d9);
or(y11, t_97, t_98);
not(z11, a9);
not(a12, b9);
not(b12, c9);
not(c12, d9);
not(t_99, t8);
not(t_100, r5);
or(d12, t_99, t_100);
not(t_101, w9);
not(t_102, s5);
or(e12, t_101, t_102);
not(t_103, q10);
not(t_104, g9);
or(f12, t_103, t_104);
not(g12, g9);
not(t_105, r10);
not(t_106, h9);
or(h12, t_105, t_106);
not(i12, h9);
not(t_107, a10);
not(t_108, v5);
or(j12, t_107, t_108);
not(t_109, b10);
not(t_110, j9);
or(k12, t_109, t_110);
not(l12, j9);
not(t_111, c10);
not(t_112, k9);
or(m12, t_111, t_112);
not(n12, k9);
not(t_113, l9);
not(t_114, o9);
or(o12, t_113, t_114);
not(t_115, m9);
not(t_116, p9);
or(p12, t_115, t_116);
not(t_117, o8);
not(t_118, a6);
or(q12, t_117, t_118);
not(r12, o9);
not(s12, p9);
not(t12, r9);
not(u12, s9);
not(v12, u9);
not(w12, v9);
not(t_119, f9);
not(t_120, j6);
or(x12, t_119, t_120);
not(t_121, i10);
not(t_122, k6);
or(y12, t_121, t_122);
not(z12, y9);
not(a13, z9);
not(t_123, i9);
not(t_124, n6);
or(b13, t_123, t_124);
not(t_125, p10);
not(t_126, r6);
or(c13, t_125, t_126);
not(t_127, o10);
not(t_128, s6);
or(d13, t_127, t_128);
not(t_129, l10);
not(t_130, t6);
or(e13, t_129, t_130);
not(t_131, g10);
not(t_132, j10);
or(f13, t_131, t_132);
not(t_133, h10);
not(t_134, k10);
or(g13, t_133, t_134);
not(t_135, x9);
not(t_136, x6);
or(h13, t_135, t_136);
not(i13, j10);
not(j13, k10);
not(t_137, f10);
not(t_138, a7);
or(k13, t_137, t_138);
not(l13, m10);
not(m13, n10);
not(t_139, e10);
not(t_140, d7);
or(n13, t_139, t_140);
not(t_141, d10);
not(t_142, f7);
or(o13, t_141, t_142);
not(t_143, t10);
not(t_144, w10);
or(p13, t_143, t_144);
not(t_145, u10);
not(t_146, x10);
or(q13, t_145, t_146);
not(r13, w10);
not(s13, x10);
not(t13, z10);
not(u13, a11);
not(t_147, q12);
not(t_148, l11);
or(v13, t_147, t_148);
not(w13, m11);
not(x13, n11);
not(t_149, q11);
not(t_150, d12);
or(y13, t_149, t_150);
not(z13, r11);
not(a14, s11);
not(t_151, b12);
not(t_152, m5);
or(b14, t_151, t_152);
not(t_153, c12);
not(t_154, n5);
or(c14, t_153, t_154);
not(t_155, x12);
not(t_156, e12);
or(d14, t_155, t_156);
not(t_157, b13);
not(t_158, j12);
or(e14, t_157, t_158);
not(t_159, r12);
not(t_160, y5);
or(f14, t_159, t_160);
not(t_161, s12);
not(t_162, z5);
or(g14, t_161, t_162);
not(t_163, h13);
not(t_164, y12);
or(h14, t_163, t_164);
not(t_165, l12);
not(t_166, o6);
or(i14, t_165, t_166);
not(t_167, n12);
not(t_168, p6);
or(j14, t_167, t_168);
not(t_169, o13);
not(t_170, c13);
or(k14, t_169, t_170);
not(t_171, n13);
not(t_172, d13);
or(l14, t_171, t_172);
not(t_173, k13);
not(t_174, e13);
or(m14, t_173, t_174);
not(t_175, i13);
not(t_176, v6);
or(n14, t_175, t_176);
not(t_177, j13);
not(t_178, w6);
or(o14, t_177, t_178);
not(t_179, g12);
not(t_180, g7);
or(p14, t_179, t_180);
not(t_181, i12);
not(t_182, h7);
or(q14, t_181, t_182);
not(t_183, r13);
not(t_184, k7);
or(r14, t_183, t_184);
not(t_185, s13);
not(t_186, l7);
or(s14, t_185, t_186);
not(t_187, t11);
not(t_188, s7);
or(t14, t_187, t_188);
not(t_189, w11);
not(t_190, t7);
or(u14, t_189, t_190);
not(v14, v13);
not(w14, y13);
not(t_191, u11);
not(t_192, t14);
or(x14, t_191, t_192);
not(t_193, v11);
not(t_194, u14);
or(y14, t_193, t_194);
not(t_195, x11);
not(t_196, b14);
or(z14, t_195, t_196);
not(t_197, y11);
not(t_198, c14);
or(a15, t_197, t_198);
not(b15, d14);
not(t_199, f12);
not(t_200, p14);
or(c15, t_199, t_200);
not(t_201, h12);
not(t_202, q14);
or(d15, t_201, t_202);
not(e15, e14);
not(t_203, k12);
not(t_204, i14);
or(f15, t_203, t_204);
not(t_205, m12);
not(t_206, j14);
or(g15, t_205, t_206);
not(t_207, o12);
not(t_208, f14);
or(h15, t_207, t_208);
not(t_209, p12);
not(t_210, g14);
or(i15, t_209, t_210);
not(t_211, q9);
not(t_212, d14);
or(j15, t_211, t_212);
not(t_213, t9);
not(t_214, y13);
or(k15, t_213, t_214);
not(l15, h14);
not(m15, k14);
not(n15, l14);
not(o15, m14);
not(t_215, f13);
not(t_216, n14);
or(p15, t_215, t_216);
not(t_217, g13);
not(t_218, o14);
or(q15, t_217, t_218);
not(t_219, s10);
not(t_220, h14);
or(r15, t_219, t_220);
not(t_221, p13);
not(t_222, r14);
or(s15, t_221, t_222);
not(t_223, q13);
not(t_224, s14);
or(t15, t_223, t_224);
not(t_225, v10);
not(t_226, m14);
or(u15, t_225, t_226);
not(t_227, y10);
not(t_228, l14);
or(v15, t_227, t_228);
not(t_229, f11);
not(t_230, c15);
or(w15, t_229, t_230);
not(t_231, g11);
not(t_232, d15);
or(x15, t_231, t_232);
not(y15, v14);
not(z15, x14);
not(a16, y14);
not(b16, z14);
not(c16, a15);
not(t_233, z11);
not(t_234, f15);
or(d16, t_233, t_234);
not(t_235, a12);
not(t_236, g15);
or(e16, t_235, t_236);
not(f16, c15);
not(g16, d15);
not(h16, e15);
not(i16, f15);
not(j16, g15);
not(k16, h15);
not(l16, i15);
not(t_237, b15);
not(t_238, d6);
or(m16, t_237, t_238);
not(t_239, t12);
not(t_240, h15);
or(n16, t_239, t_240);
not(t_241, u12);
not(t_242, i15);
or(o16, t_241, t_242);
not(t_243, w14);
not(t_244, g6);
or(p16, t_243, t_244);
not(t_245, v12);
not(t_246, z14);
or(q16, t_245, t_246);
not(t_247, w12);
not(t_248, a15);
or(r16, t_247, t_248);
buf(s16, m15);
buf(t16, m15);
not(u16, p15);
not(v16, q15);
not(t_249, l13);
not(t_250, p15);
or(w16, t_249, t_250);
not(t_251, m13);
not(t_252, q15);
or(x16, t_251, t_252);
not(t_253, l15);
not(t_254, i7);
or(y16, t_253, t_254);
not(z16, s15);
not(a17, t15);
not(t_255, o15);
not(t_256, m7);
or(b17, t_255, t_256);
not(t_257, n15);
not(t_258, p7);
or(c17, t_257, t_258);
not(t_259, t13);
not(t_260, s15);
or(d17, t_259, t_260);
not(t_261, u13);
not(t_262, t15);
or(e17, t_261, t_262);
not(t_263, f16);
not(t_264, j8);
or(f17, t_263, t_264);
not(t_265, g16);
not(t_266, k8);
or(g17, t_265, t_266);
not(h17, a16);
not(t_267, i16);
not(t_268, a9);
or(i17, t_267, t_268);
not(t_269, j16);
not(t_270, b9);
or(j17, t_269, t_270);
not(t_271, m16);
not(t_272, j15);
or(k17, t_271, t_272);
not(t_273, k16);
not(t_274, r9);
or(l17, t_273, t_274);
not(t_275, l16);
not(t_276, s9);
or(m17, t_275, t_276);
not(t_277, p16);
not(t_278, k15);
or(n17, t_277, t_278);
not(t_279, b16);
not(t_280, u9);
or(o17, t_279, t_280);
not(t_281, c16);
not(t_282, v9);
or(p17, t_281, t_282);
not(q17, s16);
not(r17, t16);
not(t_283, u16);
not(t_284, m10);
or(s17, t_283, t_284);
not(t_285, v16);
not(t_286, n10);
or(t17, t_285, t_286);
not(t_287, y16);
not(t_288, r15);
or(u17, t_287, t_288);
not(t_289, b17);
not(t_290, u15);
or(v17, t_289, t_290);
not(t_291, c17);
not(t_292, v15);
or(w17, t_291, t_292);
not(t_293, z16);
not(t_294, z10);
or(x17, t_293, t_294);
not(t_295, a17);
not(t_296, a11);
or(y17, t_295, t_296);
not(t_297, f17);
not(t_298, w15);
or(z17, t_297, t_298);
not(t_299, g17);
not(t_300, x15);
or(a18, t_299, t_300);
not(t_301, i17);
not(t_302, d16);
or(b18, t_301, t_302);
not(t_303, j17);
not(t_304, e16);
or(c18, t_303, t_304);
not(d18, k17);
not(t_305, l17);
not(t_306, n16);
or(e18, t_305, t_306);
not(t_307, m17);
not(t_308, o16);
or(f18, t_307, t_308);
not(g18, n17);
not(t_309, o17);
not(t_310, q16);
or(h18, t_309, t_310);
not(t_311, p17);
not(t_312, r16);
or(i18, t_311, t_312);
not(t_313, s17);
not(t_314, w16);
or(j18, t_313, t_314);
not(t_315, t17);
not(t_316, x16);
or(k18, t_315, t_316);
not(l18, u17);
not(m18, v17);
not(n18, w17);
not(t_317, x17);
not(t_318, d17);
or(o18, t_317, t_318);
not(t_319, y17);
not(t_320, e17);
or(p18, t_319, t_320);
not(q18, z17);
not(r18, a18);
not(t_321, g18);
not(t_322, b18);
or(s18, t_321, t_322);
not(t18, b18);
not(u18, c18);
not(t_323, m18);
not(t_324, k17);
or(v18, t_323, t_324);
not(w18, e18);
not(x18, f18);
buf(y18, h18);
buf(z18, h18);
buf(a19, h18);
not(b19, i18);
buf(c19, j18);
buf(d19, j18);
not(e19, k18);
not(f19, l18);
not(t_325, d18);
not(t_326, v17);
or(g19, t_325, t_326);
buf(h19, o18);
buf(i19, o18);
not(j19, p18);
not(k19, r18);
not(t_327, f19);
not(t_328, u18);
or(l19, t_327, t_328);
not(m19, u18);
not(t_329, v18);
not(t_330, g19);
or(n19, t_329, t_330);
buf(o19, x18);
buf(p19, x18);
buf(q19, x18);
not(t_331, t18);
not(t_332, n17);
or(r19, t_331, t_332);
not(s19, y18);
not(t19, z18);
buf(u19, a19);
buf(v19, a19);
buf(w19, b19);
buf(x19, b19);
not(t_333, z12);
not(t_334, y18);
or(y19, t_333, t_334);
not(t_335, a13);
not(t_336, z18);
or(z19, t_335, t_336);
not(a20, c19);
not(b20, d19);
buf(c20, e19);
buf(d20, e19);
not(e20, h19);
not(f20, i19);
buf(g20, j19);
buf(h20, j19);
not(t_337, r8);
not(t_338, n19);
or(i20, t_337, t_338);
not(t_339, r19);
not(t_340, s18);
or(j20, t_339, t_340);
not(k20, n19);
not(t_341, w18);
not(t_342, x19);
or(l20, t_341, t_342);
buf(m20, o19);
buf(n20, o19);
not(o20, p19);
not(p20, q19);
not(q20, u19);
not(r20, v19);
buf(s20, w19);
buf(t20, w19);
not(u20, x19);
not(t_343, s19);
not(t_344, y9);
or(v20, t_343, t_344);
not(t_345, t19);
not(t_346, z9);
or(w20, t_345, t_346);
not(t_347, a20);
not(t_348, g20);
or(x20, t_347, t_348);
not(t_349, b20);
not(t_350, h20);
or(y20, t_349, t_350);
not(z20, c20);
not(a21, d20);
not(t_351, m19);
not(t_352, l18);
or(b21, t_351, t_352);
not(c21, g20);
not(d21, h20);
not(t_353, k20);
not(t_354, j5);
or(e21, t_353, t_354);
not(f21, j20);
not(t_355, b21);
not(t_356, l19);
or(g21, t_355, t_356);
not(t_357, u20);
not(t_358, e18);
or(h21, t_357, t_358);
not(i21, m20);
not(j21, n20);
not(t_359, q20);
not(t_360, p19);
or(k21, t_359, t_360);
not(t_361, r20);
not(t_362, q19);
or(l21, t_361, t_362);
not(t_363, o20);
not(t_364, u19);
or(m21, t_363, t_364);
not(t_365, p20);
not(t_366, v19);
or(n21, t_365, t_366);
not(o21, s20);
not(p21, t20);
not(t_367, v20);
not(t_368, y19);
or(q21, t_367, t_368);
not(t_369, w20);
not(t_370, z19);
or(r21, t_369, t_370);
not(t_371, c21);
not(t_372, c19);
or(s21, t_371, t_372);
not(t_373, d21);
not(t_374, d19);
or(t21, t_373, t_374);
not(t_375, n18);
not(t_376, j20);
or(u21, t_375, t_376);
not(t_377, e20);
not(t_378, s20);
or(v21, t_377, t_378);
not(t_379, f20);
not(t_380, t20);
or(w21, t_379, t_380);
not(t_381, h11);
not(t_382, q21);
or(x21, t_381, t_382);
not(t_383, i11);
not(t_384, r21);
or(y21, t_383, t_384);
not(t_385, y15);
not(t_386, g21);
or(z21, t_385, t_386);
not(t_387, e21);
not(t_388, i20);
or(a22, t_387, t_388);
not(b22, g21);
not(t_389, h21);
not(t_390, l20);
or(c22, t_389, t_390);
not(t_391, m21);
not(t_392, k21);
or(d22, t_391, t_392);
not(t_393, n21);
not(t_394, l21);
or(e22, t_393, t_394);
not(f22, q21);
not(g22, r21);
not(t_395, s21);
not(t_396, x20);
or(h22, t_395, t_396);
not(t_397, t21);
not(t_398, y20);
or(i22, t_397, t_398);
not(t_399, f21);
not(t_400, w17);
or(j22, t_399, t_400);
not(t_401, o21);
not(t_402, h19);
or(k22, t_401, t_402);
not(t_403, p21);
not(t_404, i19);
or(l22, t_403, t_404);
not(t_405, r2);
not(t_406, a22);
or(m22, t_405, t_406);
not(t_407, f22);
not(t_408, l8);
or(n22, t_407, t_408);
not(t_409, g22);
not(t_410, m8);
or(o22, t_409, t_410);
not(t_411, b22);
not(t_412, v14);
or(p22, t_411, t_412);
buf(q22, a22);
not(t_413, h16);
not(t_414, c22);
or(r22, t_413, t_414);
not(s22, c22);
not(t22, d22);
not(u22, e22);
not(t_415, q17);
not(t_416, h22);
or(v22, t_415, t_416);
not(t_417, r17);
not(t_418, i22);
or(w22, t_417, t_418);
not(x22, h22);
not(y22, i22);
not(t_419, z20);
not(t_420, d22);
or(z22, t_419, t_420);
not(t_421, a21);
not(t_422, e22);
or(a23, t_421, t_422);
not(t_423, j22);
not(t_424, u21);
or(b23, t_423, t_424);
not(t_425, v21);
not(t_426, k22);
or(c23, t_425, t_426);
not(t_427, w21);
not(t_428, l22);
or(d23, t_427, t_428);
not(t_429, r2);
not(t_430, b23);
or(e23, t_429, t_430);
buf(f23, m22);
buf(g23, m22);
not(t_431, n22);
not(t_432, x21);
or(h23, t_431, t_432);
not(t_433, o22);
not(t_434, y21);
or(i23, t_433, t_434);
not(t_435, p22);
not(t_436, z21);
or(j23, t_435, t_436);
not(k23, q22);
not(t_437, s22);
not(t_438, e15);
or(l23, t_437, t_438);
not(t_439, i21);
not(t_440, c23);
or(m23, t_439, t_440);
not(t_441, j21);
not(t_442, d23);
or(n23, t_441, t_442);
not(t_443, x22);
not(t_444, s16);
or(o23, t_443, t_444);
not(t_445, y22);
not(t_446, t16);
or(p23, t_445, t_446);
not(t_447, t22);
not(t_448, c20);
or(q23, t_447, t_448);
not(t_449, u22);
not(t_450, d20);
or(r23, t_449, t_450);
buf(s23, b23);
not(t23, c23);
not(u23, d23);
buf(v23, e23);
buf(w23, e23);
not(x23, f23);
not(y23, g23);
not(t_451, r2);
not(t_452, j23);
or(z23, t_451, t_452);
not(t_453, b8);
not(t_454, f23);
or(a24, t_453, t_454);
not(t_455, c8);
not(t_456, g23);
or(b24, t_455, t_456);
not(c24, h23);
not(d24, i23);
buf(e24, j23);
not(t_457, l23);
not(t_458, r22);
or(f24, t_457, t_458);
not(t_459, t23);
not(t_460, m20);
or(g24, t_459, t_460);
not(t_461, u23);
not(t_462, n20);
or(h24, t_461, t_462);
not(t_463, o23);
not(t_464, v22);
or(i24, t_463, t_464);
not(t_465, p23);
not(t_466, w22);
or(j24, t_465, t_466);
not(t_467, q23);
not(t_468, z22);
or(k24, t_467, t_468);
not(t_469, r23);
not(t_470, a23);
or(l24, t_469, t_470);
not(m24, s23);
not(n24, v23);
not(o24, w23);
buf(p24, z23);
buf(q24, z23);
not(t_471, x23);
not(t_472, x4);
or(r24, t_471, t_472);
not(t_473, y23);
not(t_474, y4);
or(s24, t_473, t_474);
not(t_475, d8);
not(t_476, v23);
or(t24, t_475, t_476);
not(t_477, e8);
not(t_478, w23);
or(u24, t_477, t_478);
not(v24, d24);
not(w24, e24);
not(x24, f24);
not(t_479, g24);
not(t_480, m23);
or(y24, t_479, t_480);
not(t_481, h24);
not(t_482, n23);
or(z24, t_481, t_482);
buf(a25, i24);
buf(b25, i24);
not(c25, j24);
not(d25, k24);
not(e25, l24);
and(f25, c25, r4);
and(g25, s4, x24);
not(h25, p24);
not(i25, q24);
not(t_483, r24);
not(t_484, a24);
or(j25, t_483, t_484);
not(t_485, s24);
not(t_486, b24);
or(k25, t_485, t_486);
not(t_487, n24);
not(t_488, z4);
or(l25, t_487, t_488);
not(t_489, o24);
not(t_490, a5);
or(m25, t_489, t_490);
not(t_491, k19);
not(t_492, y24);
or(n25, t_491, t_492);
not(t_493, c24);
not(t_494, a25);
or(o25, t_493, t_494);
not(t_495, v24);
not(t_496, b25);
or(p25, t_495, t_496);
not(t_497, w13);
not(t_498, p24);
or(q25, t_497, t_498);
not(t_499, x13);
not(t_500, q24);
or(r25, t_499, t_500);
not(t_501, h17);
not(t_502, e25);
or(s25, t_501, t_502);
not(t25, y24);
not(u25, z24);
not(v25, a25);
not(w25, b25);
not(x25, e25);
not(y25, f25);
not(z25, g25);
not(a26, j25);
buf(b26, j25);
not(c26, k25);
not(t_503, l25);
not(t_504, t24);
or(d26, t_503, t_504);
not(t_505, m25);
not(t_506, u24);
or(e26, t_505, t_506);
not(t_507, q18);
not(t_508, u25);
or(f26, t_507, t_508);
not(t_509, t25);
not(t_510, r18);
or(g26, t_509, t_510);
not(t_511, v25);
not(t_512, h23);
or(h26, t_511, t_512);
not(t_513, w25);
not(t_514, d24);
or(i26, t_513, t_514);
not(t_515, h25);
not(t_516, m11);
or(j26, t_515, t_516);
not(t_517, i25);
not(t_518, n11);
or(k26, t_517, t_518);
not(t_519, x25);
not(t_520, a16);
or(l26, t_519, t_520);
not(m26, u25);
not(n26, d26);
buf(o26, d26);
not(p26, e26);
not(t_521, m26);
not(t_522, z17);
or(q26, t_521, t_522);
not(t_523, n25);
not(t_524, g26);
or(r26, t_523, t_524);
not(t_525, o25);
not(t_526, h26);
or(s26, t_525, t_526);
not(t_527, p25);
not(t_528, i26);
or(t26, t_527, t_528);
not(t_529, j26);
not(t_530, q25);
or(u26, t_529, t_530);
not(t_531, k26);
not(t_532, r25);
or(v26, t_531, t_532);
not(t_533, s25);
not(t_534, l26);
or(w26, t_533, t_534);
not(t_535, r2);
not(t_536, w26);
or(x26, t_535, t_536);
and(y26, a26, n26);
and(z26, a26, o26);
and(a27, b26, n26);
and(b27, b26, o26);
not(t_537, f26);
not(t_538, q26);
or(c27, t_537, t_538);
not(d27, r26);
not(e27, s26);
not(f27, t26);
not(g27, u26);
buf(h27, u26);
not(i27, v26);
not(t_539, r2);
not(t_540, f27);
or(j27, t_539, t_540);
not(t_541, r2);
not(t_542, c27);
or(k27, t_541, t_542);
buf(l27, x26);
buf(m27, x26);
buf(n27, j27);
buf(o27, j27);
buf(p27, k27);
buf(q27, k27);
not(r27, l27);
not(s27, m27);
not(t_543, f8);
not(t_544, l27);
or(t27, t_543, t_544);
not(t_545, g8);
not(t_546, m27);
or(u27, t_545, t_546);
not(v27, n27);
not(w27, o27);
not(x27, p27);
not(y27, q27);
not(t_547, r27);
not(t_548, b5);
or(z27, t_547, t_548);
not(t_549, s27);
not(t_550, c5);
or(a28, t_549, t_550);
not(t_551, h8);
not(t_552, p27);
or(b28, t_551, t_552);
not(t_553, i8);
not(t_554, q27);
or(c28, t_553, t_554);
not(t_555, z13);
not(t_556, n27);
or(d28, t_555, t_556);
not(t_557, a14);
not(t_558, o27);
or(e28, t_557, t_558);
not(t_559, z27);
not(t_560, t27);
or(f28, t_559, t_560);
not(t_561, a28);
not(t_562, u27);
or(g28, t_561, t_562);
not(t_563, x27);
not(t_564, d5);
or(h28, t_563, t_564);
not(t_565, y27);
not(t_566, e5);
or(i28, t_565, t_566);
not(t_567, v27);
not(t_568, r11);
or(j28, t_567, t_568);
not(t_569, w27);
not(t_570, s11);
or(k28, t_569, t_570);
not(l28, f28);
buf(m28, f28);
not(n28, g28);
not(t_571, h28);
not(t_572, b28);
or(o28, t_571, t_572);
not(t_573, i28);
not(t_574, c28);
or(p28, t_573, t_574);
not(t_575, j28);
not(t_576, d28);
or(q28, t_575, t_576);
not(t_577, k28);
not(t_578, e28);
or(r28, t_577, t_578);
not(s28, o28);
not(t28, p28);
and(u28, k11, o28);
and(v28, g27, l28);
and(w28, g27, m28);
and(x28, h27, l28);
and(y28, h27, m28);
and(z28, p11, q28);
not(a29, q28);
not(b29, r28);
and(c29, j11, s28);
and(d29, k11, s28);
buf(e29, u28);
buf(f29, u28);
not(t_579, n8);
not(t_580, b29);
not(t_581, t28);
not(t_582, s8);
not(t_583, n28);
not(t_584, p26);
not(t_585, c26);
not(t_586, i27);
or(g29, t_579, t_580, t_581, t_582, t_583, t_584, t_585, t_586);
and(h29, o11, a29);
and(i29, p11, a29);
buf(j29, z28);
buf(k29, z28);
and(l29, f2, m2, g29);
not(t_587, v7);
not(t_588, y26);
not(t_589, v28);
not(t_590, d29);
not(t_591, k29);
or(m29, t_587, t_588, t_589, t_590, t_591);
not(t_592, v7);
not(t_593, y26);
not(t_594, v28);
not(t_595, f29);
not(t_596, i29);
or(n29, t_592, t_593, t_594, t_595, t_596);
not(t_597, v7);
not(t_598, y26);
not(t_599, w28);
not(t_600, d29);
not(t_601, i29);
or(o29, t_597, t_598, t_599, t_600, t_601);
not(t_602, v7);
not(t_603, z26);
not(t_604, v28);
not(t_605, d29);
not(t_606, i29);
or(p29, t_602, t_603, t_604, t_605, t_606);
not(t_607, v7);
not(t_608, a27);
not(t_609, v28);
not(t_610, d29);
not(t_611, i29);
or(q29, t_607, t_608, t_609, t_610, t_611);
not(t_612, v7);
not(t_613, y26);
not(t_614, x28);
not(t_615, d29);
not(t_616, i29);
or(r29, t_612, t_613, t_614, t_615, t_616);
not(t_617, v7);
not(t_618, y26);
not(t_619, v28);
not(t_620, c29);
not(t_621, i29);
or(s29, t_617, t_618, t_619, t_620, t_621);
not(t_622, v7);
not(t_623, y26);
not(t_624, v28);
not(t_625, d29);
not(t_626, h29);
or(t29, t_622, t_623, t_624, t_625, t_626);
not(t_627, d11);
not(t_628, y26);
not(t_629, w28);
not(t_630, e29);
not(t_631, j29);
or(u29, t_627, t_628, t_629, t_630, t_631);
not(t_632, d11);
not(t_633, z26);
not(t_634, v28);
not(t_635, e29);
not(t_636, j29);
or(v29, t_632, t_633, t_634, t_635, t_636);
not(t_637, d11);
not(t_638, a27);
not(t_639, v28);
not(t_640, e29);
not(t_641, j29);
or(w29, t_637, t_638, t_639, t_640, t_641);
not(t_642, d11);
not(t_643, y26);
not(t_644, x28);
not(t_645, e29);
not(t_646, j29);
or(x29, t_642, t_643, t_644, t_645, t_646);
not(t_647, d11);
not(t_648, z26);
not(t_649, w28);
not(t_650, d29);
not(t_651, j29);
or(y29, t_647, t_648, t_649, t_650, t_651);
not(t_652, d11);
not(t_653, a27);
not(t_654, w28);
not(t_655, d29);
not(t_656, k29);
or(z29, t_652, t_653, t_654, t_655, t_656);
not(t_657, d11);
not(t_658, y26);
not(t_659, y28);
not(t_660, d29);
not(t_661, k29);
or(a30, t_657, t_658, t_659, t_660, t_661);
not(t_662, d11);
not(t_663, b27);
not(t_664, v28);
not(t_665, d29);
not(t_666, k29);
or(b30, t_662, t_663, t_664, t_665, t_666);
and(c30, j29, e29, w28, y26, d11);
and(d30, j29, e29, v28, z26, d11);
and(e30, j29, e29, v28, a27, d11);
and(f30, j29, e29, x28, y26, d11);
and(g30, j29, d29, w28, z26, d11);
and(h30, k29, d29, w28, a27, d11);
and(i30, k29, d29, y28, y26, d11);
and(j30, k29, d29, v28, b27, d11);
not(t_667, e11);
not(t_668, z26);
not(t_669, x28);
not(t_670, d29);
not(t_671, k29);
or(k30, t_667, t_668, t_669, t_670, t_671);
not(t_672, e11);
not(t_673, a27);
not(t_674, y28);
not(t_675, e29);
not(t_676, k29);
or(l30, t_672, t_673, t_674, t_675, t_676);
not(t_677, e11);
not(t_678, z26);
not(t_679, w28);
not(t_680, f29);
not(t_681, i29);
or(m30, t_677, t_678, t_679, t_680, t_681);
not(t_682, e11);
not(t_683, a27);
not(t_684, w28);
not(t_685, f29);
not(t_686, i29);
or(n30, t_682, t_683, t_684, t_685, t_686);
not(t_687, e11);
not(t_688, y26);
not(t_689, y28);
not(t_690, f29);
not(t_691, i29);
or(o30, t_687, t_688, t_689, t_690, t_691);
not(t_692, e11);
not(t_693, z26);
not(t_694, x28);
not(t_695, f29);
not(t_696, i29);
or(p30, t_692, t_693, t_694, t_695, t_696);
not(t_697, e11);
not(t_698, b27);
not(t_699, w28);
not(t_700, f29);
not(t_701, k29);
or(q30, t_697, t_698, t_699, t_700, t_701);
not(t_702, e11);
not(t_703, z26);
not(t_704, y28);
not(t_705, f29);
not(t_706, k29);
or(r30, t_702, t_703, t_704, t_705, t_706);
and(s30, k29, d29, x28, z26, e11);
and(t30, k29, e29, y28, a27, e11);
and(u30, i29, f29, w28, z26, e11);
and(v30, i29, f29, w28, a27, e11);
and(w30, i29, f29, y28, y26, e11);
and(x30, i29, f29, x28, z26, e11);
and(y30, k29, f29, w28, b27, e11);
and(z30, k29, f29, y28, z26, e11);
and(a31, m29, n29, o29, p29, q29, r29, s29, t29);
and(b31, u29, v29, w29, x29, y29, z29, a30, b30);
not(t_707, b30);
not(t_708, a30);
not(t_709, z29);
not(t_710, y29);
not(t_711, x29);
not(t_712, w29);
not(t_713, v29);
not(t_714, u29);
or(c31, t_707, t_708, t_709, t_710, t_711, t_712, t_713, t_714);
not(d31, c30);
not(e31, d30);
not(f31, e30);
not(g31, f30);
not(h31, g30);
not(i31, h30);
not(j31, i30);
not(k31, j30);
and(l31, k30, l30, m30, n30, o30, p30, q30, r30);
not(t_715, r30);
not(t_716, q30);
not(t_717, p30);
not(t_718, o30);
not(t_719, n30);
not(t_720, m30);
not(t_721, l30);
not(t_722, k30);
or(m31, t_715, t_716, t_717, t_718, t_719, t_720, t_721, t_722);
not(n31, s30);
not(o31, t30);
not(p31, u30);
not(q31, v30);
not(r31, w30);
not(s31, x30);
not(t31, y30);
not(u31, z30);
not(t_723, p5);
not(t_724, z30);
or(v31, t_723, t_724);
not(t_725, t5);
not(t_726, y30);
or(w31, t_725, t_726);
not(t_727, x5);
not(t_728, x30);
or(x31, t_727, t_728);
not(t_729, b6);
not(t_730, w30);
or(y31, t_729, t_730);
not(t_731, e6);
not(t_732, v30);
or(z31, t_731, t_732);
not(t_733, h6);
not(t_734, u30);
or(a32, t_733, t_734);
not(t_735, l6);
not(t_736, t30);
or(b32, t_735, t_736);
not(t_737, q6);
not(t_738, s30);
or(c32, t_737, t_738);
not(t_739, u6);
not(t_740, j30);
or(d32, t_739, t_740);
not(t_741, y6);
not(t_742, i30);
or(e32, t_741, t_742);
not(t_743, b7);
not(t_744, h30);
or(f32, t_743, t_744);
not(t_745, e7);
not(t_746, g30);
or(g32, t_745, t_746);
not(t_747, j7);
not(t_748, f30);
or(h32, t_747, t_748);
not(t_749, n7);
not(t_750, e30);
or(i32, t_749, t_750);
not(t_751, q7);
not(t_752, d30);
or(j32, t_751, t_752);
not(t_753, u7);
not(t_754, c30);
or(k32, t_753, t_754);
and(l32, b31, l31, a31);
not(t_755, l31);
not(t_756, b31);
or(m32, t_755, t_756);
and(n32, m31, k2);
and(o32, c31, l2);
not(t_757, u31);
not(t_758, g3);
or(p32, t_757, t_758);
not(t_759, t31);
not(t_760, i3);
or(q32, t_759, t_760);
not(t_761, s31);
not(t_762, k3);
or(r32, t_761, t_762);
not(t_763, r31);
not(t_764, m3);
or(s32, t_763, t_764);
not(t_765, q31);
not(t_766, o3);
or(t32, t_765, t_766);
not(t_767, p31);
not(t_768, q3);
or(u32, t_767, t_768);
not(t_769, o31);
not(t_770, s3);
or(v32, t_769, t_770);
not(t_771, n31);
not(t_772, u3);
or(w32, t_771, t_772);
not(t_773, k31);
not(t_774, w3);
or(x32, t_773, t_774);
not(t_775, j31);
not(t_776, y3);
or(y32, t_775, t_776);
not(t_777, i31);
not(t_778, a4);
or(z32, t_777, t_778);
not(t_779, h31);
not(t_780, c4);
or(a33, t_779, t_780);
not(t_781, g31);
not(t_782, e4);
or(b33, t_781, t_782);
not(t_783, f31);
not(t_784, g4);
or(c33, t_783, t_784);
not(t_785, e31);
not(t_786, i4);
or(d33, t_785, t_786);
not(t_787, d31);
not(t_788, k4);
or(e33, t_787, t_788);
not(t_789, y25);
not(t_790, o32);
or(f33, t_789, t_790);
not(t_791, z25);
not(t_792, n32);
or(g33, t_791, t_792);
not(h33, n32);
not(i33, o32);
and(j33, f2, g29, f0, l32);
and(k33, v8, s2, m32);
and(l33, q8, s2, m32);
and(m33, b0, s2, m32);
and(n33, a0, s2, m32);
and(o33, z, s2, m32);
and(p33, y, s2, m32);
not(t_793, i33);
not(t_794, f25);
or(q33, t_793, t_794);
not(t_795, h33);
not(t_796, g25);
or(r33, t_795, t_796);
not(s33, k33);
not(t33, l33);
not(u33, m33);
not(v33, n33);
not(w33, o33);
not(x33, p33);
not(t_797, d27);
not(t_798, p33);
or(y33, t_797, t_798);
not(t_799, e27);
not(t_800, k33);
or(z33, t_799, t_800);
not(t_801, w24);
not(t_802, l33);
or(a34, t_801, t_802);
not(t_803, k23);
not(t_804, m33);
or(b34, t_803, t_804);
not(t_805, d25);
not(t_806, o33);
or(c34, t_805, t_806);
not(t_807, m24);
not(t_808, n33);
or(d34, t_807, t_808);
not(t_809, q33);
not(t_810, f33);
or(e34, t_809, t_810);
not(t_811, r33);
not(t_812, g33);
or(f34, t_811, t_812);
not(t_813, x33);
not(t_814, r26);
or(g34, t_813, t_814);
not(t_815, s33);
not(t_816, s26);
or(h34, t_815, t_816);
not(t_817, t33);
not(t_818, e24);
or(i34, t_817, t_818);
not(t_819, u33);
not(t_820, q22);
or(j34, t_819, t_820);
not(t_821, w33);
not(t_822, k24);
or(k34, t_821, t_822);
not(t_823, v33);
not(t_824, s23);
or(l34, t_823, t_824);
not(m34, e34);
not(n34, f34);
not(t_825, z7);
not(t_826, e34);
or(o34, t_825, t_826);
not(t_827, a8);
not(t_828, f34);
or(p34, t_827, t_828);
not(t_829, y33);
not(t_830, g34);
or(q34, t_829, t_830);
not(t_831, z33);
not(t_832, h34);
or(r34, t_831, t_832);
not(t_833, a34);
not(t_834, i34);
or(s34, t_833, t_834);
not(t_835, b34);
not(t_836, j34);
or(t34, t_835, t_836);
not(t_837, c34);
not(t_838, k34);
or(u34, t_837, t_838);
not(t_839, d34);
not(t_840, l34);
or(v34, t_839, t_840);
not(t_841, m34);
not(t_842, t4);
or(w34, t_841, t_842);
not(t_843, n34);
not(t_844, u4);
or(x34, t_843, t_844);
not(t_845, z15);
not(t_846, u34);
or(y34, t_845, t_846);
not(z34, u34);
not(t_847, z34);
not(t_848, x14);
or(a35, t_847, t_848);
not(t_849, a35);
not(t_850, y34);
or(b35, t_849, t_850);
endmodule
module top;
	parameter in_width = 33,
		patterns = 5000,
		step = 1;
	reg [1:in_width] in_mem[1:patterns];
	integer index;

	wire i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,
		i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,
		i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,
		i30,i31,i32;

	assign {i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,
		i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,
		i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,
		i30,i31,i32} = 
		$getpattern(in_mem[index]);

	initial $monitor($time,,o0,o1,o2,o3,o4,o5,o6,o7,o8,o9,
		o10,o11,o12,o13,o14,o15,o16,o17,o18,o19,
		o20,o21,o22,o23,o24);
	initial
		begin
			$readmemb("patt.mem", in_mem);
			for(index = 1; index <= patterns; index = index + 1)
				#step;
		end

	foobar cct(o0,o1,o2,o3,o4,o5,o6,o7,o8,o9,
		o10,o11,o12,o13,o14,o15,o16,o17,o18,o19,
		o20,o21,o22,o23,o24,i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,
		i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,
		i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,
		i30,i31,i32);
endmodule