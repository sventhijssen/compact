module foobar(p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0);
input a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0;
output p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1;
not(t_0, l9);
not(t_1, a);
and(t_2, a, t_0);
and(t_3, t_1, l9);
or(p0, t_2, t_3);
not(t_4, h9);
not(t_5, b);
and(t_6, b, t_4);
and(t_7, t_5, h9);
or(q0, t_6, t_7);
not(t_8, d9);
not(t_9, c);
and(t_10, c, t_8);
and(t_11, t_9, d9);
or(r0, t_10, t_11);
not(t_12, z8);
not(t_13, d);
and(t_14, d, t_12);
and(t_15, t_13, z8);
or(s0, t_14, t_15);
not(t_16, m9);
not(t_17, e);
and(t_18, e, t_16);
and(t_19, t_17, m9);
or(t0, t_18, t_19);
not(t_20, i9);
not(t_21, f);
and(t_22, f, t_20);
and(t_23, t_21, i9);
or(u0, t_22, t_23);
not(t_24, e9);
not(t_25, g);
and(t_26, g, t_24);
and(t_27, t_25, e9);
or(v0, t_26, t_27);
not(t_28, a9);
not(t_29, h);
and(t_30, h, t_28);
and(t_31, t_29, a9);
or(w0, t_30, t_31);
not(t_32, n9);
not(t_33, i);
and(t_34, i, t_32);
and(t_35, t_33, n9);
or(x0, t_34, t_35);
not(t_36, j9);
not(t_37, j);
and(t_38, j, t_36);
and(t_39, t_37, j9);
or(y0, t_38, t_39);
not(t_40, f9);
not(t_41, k);
and(t_42, k, t_40);
and(t_43, t_41, f9);
or(z0, t_42, t_43);
not(t_44, b9);
not(t_45, l);
and(t_46, l, t_44);
and(t_47, t_45, b9);
or(a1, t_46, t_47);
not(t_48, o9);
not(t_49, m);
and(t_50, m, t_48);
and(t_51, t_49, o9);
or(b1, t_50, t_51);
not(t_52, k9);
not(t_53, n);
and(t_54, n, t_52);
and(t_55, t_53, k9);
or(c1, t_54, t_55);
not(t_56, g9);
not(t_57, o);
and(t_58, o, t_56);
and(t_59, t_57, g9);
or(d1, t_58, t_59);
not(t_60, c9);
not(t_61, p);
and(t_62, p, t_60);
and(t_63, t_61, c9);
or(e1, t_62, t_63);
not(t_64, v8);
not(t_65, q);
and(t_66, q, t_64);
and(t_67, t_65, v8);
or(f1, t_66, t_67);
not(t_68, r8);
not(t_69, r);
and(t_70, r, t_68);
and(t_71, t_69, r8);
or(g1, t_70, t_71);
not(t_72, n8);
not(t_73, s);
and(t_74, s, t_72);
and(t_75, t_73, n8);
or(h1, t_74, t_75);
not(t_76, j8);
not(t_77, t);
and(t_78, t, t_76);
and(t_79, t_77, j8);
or(i1, t_78, t_79);
not(t_80, w8);
not(t_81, u);
and(t_82, u, t_80);
and(t_83, t_81, w8);
or(j1, t_82, t_83);
not(t_84, s8);
not(t_85, v);
and(t_86, v, t_84);
and(t_87, t_85, s8);
or(k1, t_86, t_87);
not(t_88, o8);
not(t_89, w);
and(t_90, w, t_88);
and(t_91, t_89, o8);
or(l1, t_90, t_91);
not(t_92, k8);
not(t_93, x);
and(t_94, x, t_92);
and(t_95, t_93, k8);
or(m1, t_94, t_95);
not(t_96, x8);
not(t_97, y);
and(t_98, y, t_96);
and(t_99, t_97, x8);
or(n1, t_98, t_99);
not(t_100, t8);
not(t_101, z);
and(t_102, z, t_100);
and(t_103, t_101, t8);
or(o1, t_102, t_103);
not(t_104, p8);
not(t_105, a0);
and(t_106, a0, t_104);
and(t_107, t_105, p8);
or(p1, t_106, t_107);
not(t_108, l8);
not(t_109, b0);
and(t_110, b0, t_108);
and(t_111, t_109, l8);
or(q1, t_110, t_111);
not(t_112, y8);
not(t_113, c0);
and(t_114, c0, t_112);
and(t_115, t_113, y8);
or(r1, t_114, t_115);
not(t_116, u8);
not(t_117, d0);
and(t_118, d0, t_116);
and(t_119, t_117, u8);
or(s1, t_118, t_119);
not(t_120, q8);
not(t_121, e0);
and(t_122, e0, t_120);
and(t_123, t_121, q8);
or(t1, t_122, t_123);
not(t_124, m8);
not(t_125, f0);
and(t_126, f0, t_124);
and(t_127, t_125, m8);
or(u1, t_126, t_127);
and(b3, n0, o0);
and(c3, m0, o0);
and(d3, l0, o0);
and(e3, k0, o0);
and(f3, j0, o0);
and(g3, i0, o0);
and(h3, h0, o0);
and(i3, g0, o0);
not(t_128, f0);
not(t_129, e0);
and(t_130, e0, t_128);
and(t_131, t_129, f0);
or(j3, t_130, t_131);
not(t_132, d0);
not(t_133, c0);
and(t_134, c0, t_132);
and(t_135, t_133, d0);
or(k3, t_134, t_135);
not(t_136, f0);
not(t_137, b0);
and(t_138, b0, t_136);
and(t_139, t_137, f0);
or(l3, t_138, t_139);
not(t_140, e0);
not(t_141, a0);
and(t_142, a0, t_140);
and(t_143, t_141, e0);
or(m3, t_142, t_143);
not(t_144, b0);
not(t_145, a0);
and(t_146, a0, t_144);
and(t_147, t_145, b0);
or(n3, t_146, t_147);
not(t_148, d0);
not(t_149, z);
and(t_150, z, t_148);
and(t_151, t_149, d0);
or(o3, t_150, t_151);
not(t_152, c0);
not(t_153, y);
and(t_154, y, t_152);
and(t_155, t_153, c0);
or(p3, t_154, t_155);
not(t_156, z);
not(t_157, y);
and(t_158, y, t_156);
and(t_159, t_157, z);
or(q3, t_158, t_159);
not(t_160, x);
not(t_161, w);
and(t_162, w, t_160);
and(t_163, t_161, x);
or(r3, t_162, t_163);
not(t_164, v);
not(t_165, u);
and(t_166, u, t_164);
and(t_167, t_165, v);
or(s3, t_166, t_167);
not(t_168, x);
not(t_169, t);
and(t_170, t, t_168);
and(t_171, t_169, x);
or(t3, t_170, t_171);
not(t_172, w);
not(t_173, s);
and(t_174, s, t_172);
and(t_175, t_173, w);
or(u3, t_174, t_175);
not(t_176, t);
not(t_177, s);
and(t_178, s, t_176);
and(t_179, t_177, t);
or(v3, t_178, t_179);
not(t_180, v);
not(t_181, r);
and(t_182, r, t_180);
and(t_183, t_181, v);
or(w3, t_182, t_183);
not(t_184, u);
not(t_185, q);
and(t_186, q, t_184);
and(t_187, t_185, u);
or(x3, t_186, t_187);
not(t_188, r);
not(t_189, q);
and(t_190, q, t_188);
and(t_191, t_189, r);
or(y3, t_190, t_191);
not(t_192, p);
not(t_193, o);
and(t_194, o, t_192);
and(t_195, t_193, p);
or(z3, t_194, t_195);
not(t_196, n);
not(t_197, m);
and(t_198, m, t_196);
and(t_199, t_197, n);
or(a4, t_198, t_199);
not(t_200, p);
not(t_201, l);
and(t_202, l, t_200);
and(t_203, t_201, p);
or(b4, t_202, t_203);
not(t_204, o);
not(t_205, k);
and(t_206, k, t_204);
and(t_207, t_205, o);
or(c4, t_206, t_207);
not(t_208, l);
not(t_209, k);
and(t_210, k, t_208);
and(t_211, t_209, l);
or(d4, t_210, t_211);
not(t_212, n);
not(t_213, j);
and(t_214, j, t_212);
and(t_215, t_213, n);
or(e4, t_214, t_215);
not(t_216, m);
not(t_217, i);
and(t_218, i, t_216);
and(t_219, t_217, m);
or(f4, t_218, t_219);
not(t_220, j);
not(t_221, i);
and(t_222, i, t_220);
and(t_223, t_221, j);
or(g4, t_222, t_223);
not(t_224, h);
not(t_225, g);
and(t_226, g, t_224);
and(t_227, t_225, h);
or(h4, t_226, t_227);
not(t_228, f);
not(t_229, e);
and(t_230, e, t_228);
and(t_231, t_229, f);
or(i4, t_230, t_231);
not(t_232, h);
not(t_233, d);
and(t_234, d, t_232);
and(t_235, t_233, h);
or(j4, t_234, t_235);
not(t_236, g);
not(t_237, c);
and(t_238, c, t_236);
and(t_239, t_237, g);
or(k4, t_238, t_239);
not(t_240, d);
not(t_241, c);
and(t_242, c, t_240);
and(t_243, t_241, d);
or(l4, t_242, t_243);
not(t_244, f);
not(t_245, b);
and(t_246, b, t_244);
and(t_247, t_245, f);
or(m4, t_246, t_247);
not(t_248, e);
not(t_249, a);
and(t_250, a, t_248);
and(t_251, t_249, e);
or(n4, t_250, t_251);
not(t_252, b);
not(t_253, a);
and(t_254, a, t_252);
and(t_255, t_253, b);
or(o4, t_254, t_255);
not(t_256, j3);
not(t_257, k3);
and(t_258, k3, t_256);
and(t_259, t_257, j3);
or(p4, t_258, t_259);
not(t_260, l3);
not(t_261, t3);
and(t_262, t3, t_260);
and(t_263, t_261, l3);
or(q4, t_262, t_263);
not(t_264, m3);
not(t_265, u3);
and(t_266, u3, t_264);
and(t_267, t_265, m3);
or(r4, t_266, t_267);
not(t_268, n3);
not(t_269, q3);
and(t_270, q3, t_268);
and(t_271, t_269, n3);
or(s4, t_270, t_271);
not(t_272, o3);
not(t_273, w3);
and(t_274, w3, t_272);
and(t_275, t_273, o3);
or(t4, t_274, t_275);
not(t_276, p3);
not(t_277, x3);
and(t_278, x3, t_276);
and(t_279, t_277, p3);
or(u4, t_278, t_279);
not(t_280, r3);
not(t_281, s3);
and(t_282, s3, t_280);
and(t_283, t_281, r3);
or(v4, t_282, t_283);
not(t_284, v3);
not(t_285, y3);
and(t_286, y3, t_284);
and(t_287, t_285, v3);
or(w4, t_286, t_287);
not(t_288, z3);
not(t_289, a4);
and(t_290, a4, t_288);
and(t_291, t_289, z3);
or(x4, t_290, t_291);
not(t_292, b4);
not(t_293, j4);
and(t_294, j4, t_292);
and(t_295, t_293, b4);
or(y4, t_294, t_295);
not(t_296, c4);
not(t_297, k4);
and(t_298, k4, t_296);
and(t_299, t_297, c4);
or(z4, t_298, t_299);
not(t_300, d4);
not(t_301, g4);
and(t_302, g4, t_300);
and(t_303, t_301, d4);
or(a5, t_302, t_303);
not(t_304, e4);
not(t_305, m4);
and(t_306, m4, t_304);
and(t_307, t_305, e4);
or(b5, t_306, t_307);
not(t_308, f4);
not(t_309, n4);
and(t_310, n4, t_308);
and(t_311, t_309, f4);
or(c5, t_310, t_311);
not(t_312, h4);
not(t_313, i4);
and(t_314, i4, t_312);
and(t_315, t_313, h4);
or(d5, t_314, t_315);
not(t_316, l4);
not(t_317, o4);
and(t_318, o4, t_316);
and(t_319, t_317, l4);
or(e5, t_318, t_319);
not(t_320, p4);
not(t_321, s4);
and(t_322, s4, t_320);
and(t_323, t_321, p4);
or(f5, t_322, t_323);
not(t_324, p4);
not(t_325, v4);
and(t_326, v4, t_324);
and(t_327, t_325, p4);
or(g5, t_326, t_327);
not(t_328, s4);
not(t_329, w4);
and(t_330, w4, t_328);
and(t_331, t_329, s4);
or(h5, t_330, t_331);
not(t_332, v4);
not(t_333, w4);
and(t_334, w4, t_332);
and(t_335, t_333, v4);
or(i5, t_334, t_335);
not(t_336, x4);
not(t_337, a5);
and(t_338, a5, t_336);
and(t_339, t_337, x4);
or(j5, t_338, t_339);
not(t_340, x4);
not(t_341, d5);
and(t_342, d5, t_340);
and(t_343, t_341, x4);
or(k5, t_342, t_343);
not(t_344, a5);
not(t_345, e5);
and(t_346, e5, t_344);
and(t_347, t_345, a5);
or(l5, t_346, t_347);
not(t_348, d5);
not(t_349, e5);
and(t_350, e5, t_348);
and(t_351, t_349, d5);
or(m5, t_350, t_351);
not(t_352, k5);
not(t_353, b3);
and(t_354, b3, t_352);
and(t_355, t_353, k5);
or(n5, t_354, t_355);
not(t_356, l5);
not(t_357, c3);
and(t_358, c3, t_356);
and(t_359, t_357, l5);
or(o5, t_358, t_359);
not(t_360, j5);
not(t_361, d3);
and(t_362, d3, t_360);
and(t_363, t_361, j5);
or(p5, t_362, t_363);
not(t_364, m5);
not(t_365, e3);
and(t_366, e3, t_364);
and(t_367, t_365, m5);
or(q5, t_366, t_367);
not(t_368, g5);
not(t_369, f3);
and(t_370, f3, t_368);
and(t_371, t_369, g5);
or(r5, t_370, t_371);
not(t_372, h5);
not(t_373, g3);
and(t_374, g3, t_372);
and(t_375, t_373, h5);
or(s5, t_374, t_375);
not(t_376, f5);
not(t_377, h3);
and(t_378, h3, t_376);
and(t_379, t_377, f5);
or(t5, t_378, t_379);
not(t_380, i5);
not(t_381, i3);
and(t_382, i3, t_380);
and(t_383, t_381, i5);
or(u5, t_382, t_383);
not(t_384, n5);
not(t_385, q4);
and(t_386, q4, t_384);
and(t_387, t_385, n5);
or(v5, t_386, t_387);
not(t_388, o5);
not(t_389, r4);
and(t_390, r4, t_388);
and(t_391, t_389, o5);
or(w5, t_390, t_391);
not(t_392, p5);
not(t_393, t4);
and(t_394, t4, t_392);
and(t_395, t_393, p5);
or(x5, t_394, t_395);
not(t_396, q5);
not(t_397, u4);
and(t_398, u4, t_396);
and(t_399, t_397, q5);
or(y5, t_398, t_399);
not(t_400, r5);
not(t_401, y4);
and(t_402, y4, t_400);
and(t_403, t_401, r5);
or(z5, t_402, t_403);
not(t_404, s5);
not(t_405, z4);
and(t_406, z4, t_404);
and(t_407, t_405, s5);
or(a6, t_406, t_407);
not(t_408, t5);
not(t_409, b5);
and(t_410, b5, t_408);
and(t_411, t_409, t5);
or(b6, t_410, t_411);
not(t_412, u5);
not(t_413, c5);
and(t_414, c5, t_412);
and(t_415, t_413, u5);
or(c6, t_414, t_415);
not(d6, v5);
not(e6, v5);
not(f6, v5);
not(g6, v5);
not(h6, v5);
not(i6, w5);
not(j6, w5);
not(k6, w5);
not(l6, w5);
not(m6, w5);
not(n6, x5);
not(o6, x5);
not(p6, x5);
not(q6, x5);
not(r6, x5);
not(s6, y5);
not(t6, y5);
not(u6, y5);
not(v6, y5);
not(w6, y5);
not(x6, z5);
not(y6, z5);
not(z6, z5);
not(a7, z5);
not(b7, z5);
not(c7, a6);
not(d7, a6);
not(e7, a6);
not(f7, a6);
not(g7, a6);
not(h7, b6);
not(i7, b6);
not(j7, b6);
not(k7, b6);
not(l7, b6);
not(m7, c6);
not(n7, c6);
not(o7, c6);
not(p7, c6);
not(q7, c6);
and(r7, s6, n6, i6, v5);
and(s7, t6, o6, w5, d6);
and(t7, u6, x5, j6, e6);
and(u7, y5, p6, k6, f6);
and(v7, m7, h7, c7, z5);
and(w7, n7, i7, a6, x6);
and(x7, o7, b6, d7, y6);
and(y7, c6, j7, e7, z6);
or(z7, u7, t7, s7, r7);
or(a8, y7, x7, w7, v7);
and(b8, y5, r6, l6, v5, a8);
and(c8, w6, x5, m6, v5, a8);
and(d8, y5, q6, w5, g6, a8);
and(e8, v6, x5, w5, h6, a8);
and(f8, c6, l7, f7, z5, z7);
and(g8, q7, b6, g7, z5, z7);
and(h8, c6, k7, a6, a7, z7);
and(i8, p7, b6, a6, b7, z7);
and(j8, v5, h8);
and(k8, v5, f8);
and(l8, v5, i8);
and(m8, v5, g8);
and(n8, w5, h8);
and(o8, w5, f8);
and(p8, w5, i8);
and(q8, w5, g8);
and(r8, x5, h8);
and(s8, x5, f8);
and(t8, x5, i8);
and(u8, x5, g8);
and(v8, y5, h8);
and(w8, y5, f8);
and(x8, y5, i8);
and(y8, y5, g8);
and(z8, z5, d8);
and(a9, z5, b8);
and(b9, z5, e8);
and(c9, z5, c8);
and(d9, a6, d8);
and(e9, a6, b8);
and(f9, a6, e8);
and(g9, a6, c8);
and(h9, b6, d8);
and(i9, b6, b8);
and(j9, b6, e8);
and(k9, b6, c8);
and(l9, c6, d8);
and(m9, c6, b8);
and(n9, c6, e8);
and(o9, c6, c8);
endmodule
module top;
	parameter in_width = 41,
		patterns = 5000,
		step = 1;
	reg [1:in_width] in_mem[1:patterns];
	integer index;

	wire i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,
		i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,
		i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,
		i30,i31,i32,i33,i34,i35,i36,i37,i38,i39,
		i40;

	assign {i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,
		i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,
		i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,
		i30,i31,i32,i33,i34,i35,i36,i37,i38,i39,
		i40} = 
		$getpattern(in_mem[index]);

	initial $monitor($time,,o0,o1,o2,o3,o4,o5,o6,o7,o8,o9,
		o10,o11,o12,o13,o14,o15,o16,o17,o18,o19,
		o20,o21,o22,o23,o24,o25,o26,o27,o28,o29,
		o30,o31);
	initial
		begin
			$readmemb("patt.mem", in_mem);
			for(index = 1; index <= patterns; index = index + 1)
				#step;
		end

	foobar cct(o0,o1,o2,o3,o4,o5,o6,o7,o8,o9,
		o10,o11,o12,o13,o14,o15,o16,o17,o18,o19,
		o20,o21,o22,o23,o24,o25,o26,o27,o28,o29,
		o30,o31,i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,
		i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,
		i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,
		i30,i31,i32,i33,i34,i35,i36,i37,i38,i39,
		i40);
endmodule